library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sqrtROM is
    port (
        Clk    : in  std_logic;                       -- Clock signal
        en     : in  std_logic;
        Addr   : in  std_logic_vector(17 downto 0);   -- 18-bit Address input
        SqRoot : out std_logic_vector(8 downto 0);     -- 9-bit Square Root output
        data_valid : out std_logic 
    );
end entity;

architecture Behavioral of sqrtROM is
    -- ROM content: 1024 x 9-bit memory for storing square roots
    type rom_type is array (0 to 8191) of std_logic_vector(8 downto 0);

    -- Initialize ROM with precomputed square roots (truncated to 9 bits)
    constant ROM : rom_type := (
"000000000",  -- sqrt(   0) = 0
"000000001",  -- sqrt(   1) = 1
"000000001",  -- sqrt(   2) = 1
"000000010",  -- sqrt(   3) = 2
"000000010",  -- sqrt(   4) = 2
"000000010",  -- sqrt(   5) = 2
"000000010",  -- sqrt(   6) = 2
"000000011",  -- sqrt(   7) = 3
"000000011",  -- sqrt(   8) = 3
"000000011",  -- sqrt(   9) = 3
"000000011",  -- sqrt(  10) = 3
"000000011",  -- sqrt(  11) = 3
"000000011",  -- sqrt(  12) = 3
"000000100",  -- sqrt(  13) = 4
"000000100",  -- sqrt(  14) = 4
"000000100",  -- sqrt(  15) = 4
"000000100",  -- sqrt(  16) = 4
"000000100",  -- sqrt(  17) = 4
"000000100",  -- sqrt(  18) = 4
"000000100",  -- sqrt(  19) = 4
"000000100",  -- sqrt(  20) = 4
"000000101",  -- sqrt(  21) = 5
"000000101",  -- sqrt(  22) = 5
"000000101",  -- sqrt(  23) = 5
"000000101",  -- sqrt(  24) = 5
"000000101",  -- sqrt(  25) = 5
"000000101",  -- sqrt(  26) = 5
"000000101",  -- sqrt(  27) = 5
"000000101",  -- sqrt(  28) = 5
"000000101",  -- sqrt(  29) = 5
"000000101",  -- sqrt(  30) = 5
"000000110",  -- sqrt(  31) = 6
"000000110",  -- sqrt(  32) = 6
"000000110",  -- sqrt(  33) = 6
"000000110",  -- sqrt(  34) = 6
"000000110",  -- sqrt(  35) = 6
"000000110",  -- sqrt(  36) = 6
"000000110",  -- sqrt(  37) = 6
"000000110",  -- sqrt(  38) = 6
"000000110",  -- sqrt(  39) = 6
"000000110",  -- sqrt(  40) = 6
"000000110",  -- sqrt(  41) = 6
"000000110",  -- sqrt(  42) = 6
"000000111",  -- sqrt(  43) = 7
"000000111",  -- sqrt(  44) = 7
"000000111",  -- sqrt(  45) = 7
"000000111",  -- sqrt(  46) = 7
"000000111",  -- sqrt(  47) = 7
"000000111",  -- sqrt(  48) = 7
"000000111",  -- sqrt(  49) = 7
"000000111",  -- sqrt(  50) = 7
"000000111",  -- sqrt(  51) = 7
"000000111",  -- sqrt(  52) = 7
"000000111",  -- sqrt(  53) = 7
"000000111",  -- sqrt(  54) = 7
"000000111",  -- sqrt(  55) = 7
"000000111",  -- sqrt(  56) = 7
"000001000",  -- sqrt(  57) = 8
"000001000",  -- sqrt(  58) = 8
"000001000",  -- sqrt(  59) = 8
"000001000",  -- sqrt(  60) = 8
"000001000",  -- sqrt(  61) = 8
"000001000",  -- sqrt(  62) = 8
"000001000",  -- sqrt(  63) = 8
"000001000",  -- sqrt(  64) = 8
"000001000",  -- sqrt(  65) = 8
"000001000",  -- sqrt(  66) = 8
"000001000",  -- sqrt(  67) = 8
"000001000",  -- sqrt(  68) = 8
"000001000",  -- sqrt(  69) = 8
"000001000",  -- sqrt(  70) = 8
"000001000",  -- sqrt(  71) = 8
"000001000",  -- sqrt(  72) = 8
"000001001",  -- sqrt(  73) = 9
"000001001",  -- sqrt(  74) = 9
"000001001",  -- sqrt(  75) = 9
"000001001",  -- sqrt(  76) = 9
"000001001",  -- sqrt(  77) = 9
"000001001",  -- sqrt(  78) = 9
"000001001",  -- sqrt(  79) = 9
"000001001",  -- sqrt(  80) = 9
"000001001",  -- sqrt(  81) = 9
"000001001",  -- sqrt(  82) = 9
"000001001",  -- sqrt(  83) = 9
"000001001",  -- sqrt(  84) = 9
"000001001",  -- sqrt(  85) = 9
"000001001",  -- sqrt(  86) = 9
"000001001",  -- sqrt(  87) = 9
"000001001",  -- sqrt(  88) = 9
"000001001",  -- sqrt(  89) = 9
"000001001",  -- sqrt(  90) = 9
"000001010",  -- sqrt(  91) = 10
"000001010",  -- sqrt(  92) = 10
"000001010",  -- sqrt(  93) = 10
"000001010",  -- sqrt(  94) = 10
"000001010",  -- sqrt(  95) = 10
"000001010",  -- sqrt(  96) = 10
"000001010",  -- sqrt(  97) = 10
"000001010",  -- sqrt(  98) = 10
"000001010",  -- sqrt(  99) = 10
"000001010",  -- sqrt( 100) = 10
"000001010",  -- sqrt( 101) = 10
"000001010",  -- sqrt( 102) = 10
"000001010",  -- sqrt( 103) = 10
"000001010",  -- sqrt( 104) = 10
"000001010",  -- sqrt( 105) = 10
"000001010",  -- sqrt( 106) = 10
"000001010",  -- sqrt( 107) = 10
"000001010",  -- sqrt( 108) = 10
"000001010",  -- sqrt( 109) = 10
"000001010",  -- sqrt( 110) = 10
"000001011",  -- sqrt( 111) = 11
"000001011",  -- sqrt( 112) = 11
"000001011",  -- sqrt( 113) = 11
"000001011",  -- sqrt( 114) = 11
"000001011",  -- sqrt( 115) = 11
"000001011",  -- sqrt( 116) = 11
"000001011",  -- sqrt( 117) = 11
"000001011",  -- sqrt( 118) = 11
"000001011",  -- sqrt( 119) = 11
"000001011",  -- sqrt( 120) = 11
"000001011",  -- sqrt( 121) = 11
"000001011",  -- sqrt( 122) = 11
"000001011",  -- sqrt( 123) = 11
"000001011",  -- sqrt( 124) = 11
"000001011",  -- sqrt( 125) = 11
"000001011",  -- sqrt( 126) = 11
"000001011",  -- sqrt( 127) = 11
"000001011",  -- sqrt( 128) = 11
"000001011",  -- sqrt( 129) = 11
"000001011",  -- sqrt( 130) = 11
"000001011",  -- sqrt( 131) = 11
"000001011",  -- sqrt( 132) = 11
"000001100",  -- sqrt( 133) = 12
"000001100",  -- sqrt( 134) = 12
"000001100",  -- sqrt( 135) = 12
"000001100",  -- sqrt( 136) = 12
"000001100",  -- sqrt( 137) = 12
"000001100",  -- sqrt( 138) = 12
"000001100",  -- sqrt( 139) = 12
"000001100",  -- sqrt( 140) = 12
"000001100",  -- sqrt( 141) = 12
"000001100",  -- sqrt( 142) = 12
"000001100",  -- sqrt( 143) = 12
"000001100",  -- sqrt( 144) = 12
"000001100",  -- sqrt( 145) = 12
"000001100",  -- sqrt( 146) = 12
"000001100",  -- sqrt( 147) = 12
"000001100",  -- sqrt( 148) = 12
"000001100",  -- sqrt( 149) = 12
"000001100",  -- sqrt( 150) = 12
"000001100",  -- sqrt( 151) = 12
"000001100",  -- sqrt( 152) = 12
"000001100",  -- sqrt( 153) = 12
"000001100",  -- sqrt( 154) = 12
"000001100",  -- sqrt( 155) = 12
"000001100",  -- sqrt( 156) = 12
"000001101",  -- sqrt( 157) = 13
"000001101",  -- sqrt( 158) = 13
"000001101",  -- sqrt( 159) = 13
"000001101",  -- sqrt( 160) = 13
"000001101",  -- sqrt( 161) = 13
"000001101",  -- sqrt( 162) = 13
"000001101",  -- sqrt( 163) = 13
"000001101",  -- sqrt( 164) = 13
"000001101",  -- sqrt( 165) = 13
"000001101",  -- sqrt( 166) = 13
"000001101",  -- sqrt( 167) = 13
"000001101",  -- sqrt( 168) = 13
"000001101",  -- sqrt( 169) = 13
"000001101",  -- sqrt( 170) = 13
"000001101",  -- sqrt( 171) = 13
"000001101",  -- sqrt( 172) = 13
"000001101",  -- sqrt( 173) = 13
"000001101",  -- sqrt( 174) = 13
"000001101",  -- sqrt( 175) = 13
"000001101",  -- sqrt( 176) = 13
"000001101",  -- sqrt( 177) = 13
"000001101",  -- sqrt( 178) = 13
"000001101",  -- sqrt( 179) = 13
"000001101",  -- sqrt( 180) = 13
"000001101",  -- sqrt( 181) = 13
"000001101",  -- sqrt( 182) = 13
"000001110",  -- sqrt( 183) = 14
"000001110",  -- sqrt( 184) = 14
"000001110",  -- sqrt( 185) = 14
"000001110",  -- sqrt( 186) = 14
"000001110",  -- sqrt( 187) = 14
"000001110",  -- sqrt( 188) = 14
"000001110",  -- sqrt( 189) = 14
"000001110",  -- sqrt( 190) = 14
"000001110",  -- sqrt( 191) = 14
"000001110",  -- sqrt( 192) = 14
"000001110",  -- sqrt( 193) = 14
"000001110",  -- sqrt( 194) = 14
"000001110",  -- sqrt( 195) = 14
"000001110",  -- sqrt( 196) = 14
"000001110",  -- sqrt( 197) = 14
"000001110",  -- sqrt( 198) = 14
"000001110",  -- sqrt( 199) = 14
"000001110",  -- sqrt( 200) = 14
"000001110",  -- sqrt( 201) = 14
"000001110",  -- sqrt( 202) = 14
"000001110",  -- sqrt( 203) = 14
"000001110",  -- sqrt( 204) = 14
"000001110",  -- sqrt( 205) = 14
"000001110",  -- sqrt( 206) = 14
"000001110",  -- sqrt( 207) = 14
"000001110",  -- sqrt( 208) = 14
"000001110",  -- sqrt( 209) = 14
"000001110",  -- sqrt( 210) = 14
"000001111",  -- sqrt( 211) = 15
"000001111",  -- sqrt( 212) = 15
"000001111",  -- sqrt( 213) = 15
"000001111",  -- sqrt( 214) = 15
"000001111",  -- sqrt( 215) = 15
"000001111",  -- sqrt( 216) = 15
"000001111",  -- sqrt( 217) = 15
"000001111",  -- sqrt( 218) = 15
"000001111",  -- sqrt( 219) = 15
"000001111",  -- sqrt( 220) = 15
"000001111",  -- sqrt( 221) = 15
"000001111",  -- sqrt( 222) = 15
"000001111",  -- sqrt( 223) = 15
"000001111",  -- sqrt( 224) = 15
"000001111",  -- sqrt( 225) = 15
"000001111",  -- sqrt( 226) = 15
"000001111",  -- sqrt( 227) = 15
"000001111",  -- sqrt( 228) = 15
"000001111",  -- sqrt( 229) = 15
"000001111",  -- sqrt( 230) = 15
"000001111",  -- sqrt( 231) = 15
"000001111",  -- sqrt( 232) = 15
"000001111",  -- sqrt( 233) = 15
"000001111",  -- sqrt( 234) = 15
"000001111",  -- sqrt( 235) = 15
"000001111",  -- sqrt( 236) = 15
"000001111",  -- sqrt( 237) = 15
"000001111",  -- sqrt( 238) = 15
"000001111",  -- sqrt( 239) = 15
"000001111",  -- sqrt( 240) = 15
"000010000",  -- sqrt( 241) = 16
"000010000",  -- sqrt( 242) = 16
"000010000",  -- sqrt( 243) = 16
"000010000",  -- sqrt( 244) = 16
"000010000",  -- sqrt( 245) = 16
"000010000",  -- sqrt( 246) = 16
"000010000",  -- sqrt( 247) = 16
"000010000",  -- sqrt( 248) = 16
"000010000",  -- sqrt( 249) = 16
"000010000",  -- sqrt( 250) = 16
"000010000",  -- sqrt( 251) = 16
"000010000",  -- sqrt( 252) = 16
"000010000",  -- sqrt( 253) = 16
"000010000",  -- sqrt( 254) = 16
"000010000",  -- sqrt( 255) = 16
"000010000",  -- sqrt( 256) = 16
"000010000",  -- sqrt( 257) = 16
"000010000",  -- sqrt( 258) = 16
"000010000",  -- sqrt( 259) = 16
"000010000",  -- sqrt( 260) = 16
"000010000",  -- sqrt( 261) = 16
"000010000",  -- sqrt( 262) = 16
"000010000",  -- sqrt( 263) = 16
"000010000",  -- sqrt( 264) = 16
"000010000",  -- sqrt( 265) = 16
"000010000",  -- sqrt( 266) = 16
"000010000",  -- sqrt( 267) = 16
"000010000",  -- sqrt( 268) = 16
"000010000",  -- sqrt( 269) = 16
"000010000",  -- sqrt( 270) = 16
"000010000",  -- sqrt( 271) = 16
"000010000",  -- sqrt( 272) = 16
"000010001",  -- sqrt( 273) = 17
"000010001",  -- sqrt( 274) = 17
"000010001",  -- sqrt( 275) = 17
"000010001",  -- sqrt( 276) = 17
"000010001",  -- sqrt( 277) = 17
"000010001",  -- sqrt( 278) = 17
"000010001",  -- sqrt( 279) = 17
"000010001",  -- sqrt( 280) = 17
"000010001",  -- sqrt( 281) = 17
"000010001",  -- sqrt( 282) = 17
"000010001",  -- sqrt( 283) = 17
"000010001",  -- sqrt( 284) = 17
"000010001",  -- sqrt( 285) = 17
"000010001",  -- sqrt( 286) = 17
"000010001",  -- sqrt( 287) = 17
"000010001",  -- sqrt( 288) = 17
"000010001",  -- sqrt( 289) = 17
"000010001",  -- sqrt( 290) = 17
"000010001",  -- sqrt( 291) = 17
"000010001",  -- sqrt( 292) = 17
"000010001",  -- sqrt( 293) = 17
"000010001",  -- sqrt( 294) = 17
"000010001",  -- sqrt( 295) = 17
"000010001",  -- sqrt( 296) = 17
"000010001",  -- sqrt( 297) = 17
"000010001",  -- sqrt( 298) = 17
"000010001",  -- sqrt( 299) = 17
"000010001",  -- sqrt( 300) = 17
"000010001",  -- sqrt( 301) = 17
"000010001",  -- sqrt( 302) = 17
"000010001",  -- sqrt( 303) = 17
"000010001",  -- sqrt( 304) = 17
"000010001",  -- sqrt( 305) = 17
"000010001",  -- sqrt( 306) = 17
"000010010",  -- sqrt( 307) = 18
"000010010",  -- sqrt( 308) = 18
"000010010",  -- sqrt( 309) = 18
"000010010",  -- sqrt( 310) = 18
"000010010",  -- sqrt( 311) = 18
"000010010",  -- sqrt( 312) = 18
"000010010",  -- sqrt( 313) = 18
"000010010",  -- sqrt( 314) = 18
"000010010",  -- sqrt( 315) = 18
"000010010",  -- sqrt( 316) = 18
"000010010",  -- sqrt( 317) = 18
"000010010",  -- sqrt( 318) = 18
"000010010",  -- sqrt( 319) = 18
"000010010",  -- sqrt( 320) = 18
"000010010",  -- sqrt( 321) = 18
"000010010",  -- sqrt( 322) = 18
"000010010",  -- sqrt( 323) = 18
"000010010",  -- sqrt( 324) = 18
"000010010",  -- sqrt( 325) = 18
"000010010",  -- sqrt( 326) = 18
"000010010",  -- sqrt( 327) = 18
"000010010",  -- sqrt( 328) = 18
"000010010",  -- sqrt( 329) = 18
"000010010",  -- sqrt( 330) = 18
"000010010",  -- sqrt( 331) = 18
"000010010",  -- sqrt( 332) = 18
"000010010",  -- sqrt( 333) = 18
"000010010",  -- sqrt( 334) = 18
"000010010",  -- sqrt( 335) = 18
"000010010",  -- sqrt( 336) = 18
"000010010",  -- sqrt( 337) = 18
"000010010",  -- sqrt( 338) = 18
"000010010",  -- sqrt( 339) = 18
"000010010",  -- sqrt( 340) = 18
"000010010",  -- sqrt( 341) = 18
"000010010",  -- sqrt( 342) = 18
"000010011",  -- sqrt( 343) = 19
"000010011",  -- sqrt( 344) = 19
"000010011",  -- sqrt( 345) = 19
"000010011",  -- sqrt( 346) = 19
"000010011",  -- sqrt( 347) = 19
"000010011",  -- sqrt( 348) = 19
"000010011",  -- sqrt( 349) = 19
"000010011",  -- sqrt( 350) = 19
"000010011",  -- sqrt( 351) = 19
"000010011",  -- sqrt( 352) = 19
"000010011",  -- sqrt( 353) = 19
"000010011",  -- sqrt( 354) = 19
"000010011",  -- sqrt( 355) = 19
"000010011",  -- sqrt( 356) = 19
"000010011",  -- sqrt( 357) = 19
"000010011",  -- sqrt( 358) = 19
"000010011",  -- sqrt( 359) = 19
"000010011",  -- sqrt( 360) = 19
"000010011",  -- sqrt( 361) = 19
"000010011",  -- sqrt( 362) = 19
"000010011",  -- sqrt( 363) = 19
"000010011",  -- sqrt( 364) = 19
"000010011",  -- sqrt( 365) = 19
"000010011",  -- sqrt( 366) = 19
"000010011",  -- sqrt( 367) = 19
"000010011",  -- sqrt( 368) = 19
"000010011",  -- sqrt( 369) = 19
"000010011",  -- sqrt( 370) = 19
"000010011",  -- sqrt( 371) = 19
"000010011",  -- sqrt( 372) = 19
"000010011",  -- sqrt( 373) = 19
"000010011",  -- sqrt( 374) = 19
"000010011",  -- sqrt( 375) = 19
"000010011",  -- sqrt( 376) = 19
"000010011",  -- sqrt( 377) = 19
"000010011",  -- sqrt( 378) = 19
"000010011",  -- sqrt( 379) = 19
"000010011",  -- sqrt( 380) = 19
"000010100",  -- sqrt( 381) = 20
"000010100",  -- sqrt( 382) = 20
"000010100",  -- sqrt( 383) = 20
"000010100",  -- sqrt( 384) = 20
"000010100",  -- sqrt( 385) = 20
"000010100",  -- sqrt( 386) = 20
"000010100",  -- sqrt( 387) = 20
"000010100",  -- sqrt( 388) = 20
"000010100",  -- sqrt( 389) = 20
"000010100",  -- sqrt( 390) = 20
"000010100",  -- sqrt( 391) = 20
"000010100",  -- sqrt( 392) = 20
"000010100",  -- sqrt( 393) = 20
"000010100",  -- sqrt( 394) = 20
"000010100",  -- sqrt( 395) = 20
"000010100",  -- sqrt( 396) = 20
"000010100",  -- sqrt( 397) = 20
"000010100",  -- sqrt( 398) = 20
"000010100",  -- sqrt( 399) = 20
"000010100",  -- sqrt( 400) = 20
"000010100",  -- sqrt( 401) = 20
"000010100",  -- sqrt( 402) = 20
"000010100",  -- sqrt( 403) = 20
"000010100",  -- sqrt( 404) = 20
"000010100",  -- sqrt( 405) = 20
"000010100",  -- sqrt( 406) = 20
"000010100",  -- sqrt( 407) = 20
"000010100",  -- sqrt( 408) = 20
"000010100",  -- sqrt( 409) = 20
"000010100",  -- sqrt( 410) = 20
"000010100",  -- sqrt( 411) = 20
"000010100",  -- sqrt( 412) = 20
"000010100",  -- sqrt( 413) = 20
"000010100",  -- sqrt( 414) = 20
"000010100",  -- sqrt( 415) = 20
"000010100",  -- sqrt( 416) = 20
"000010100",  -- sqrt( 417) = 20
"000010100",  -- sqrt( 418) = 20
"000010100",  -- sqrt( 419) = 20
"000010100",  -- sqrt( 420) = 20
"000010101",  -- sqrt( 421) = 21
"000010101",  -- sqrt( 422) = 21
"000010101",  -- sqrt( 423) = 21
"000010101",  -- sqrt( 424) = 21
"000010101",  -- sqrt( 425) = 21
"000010101",  -- sqrt( 426) = 21
"000010101",  -- sqrt( 427) = 21
"000010101",  -- sqrt( 428) = 21
"000010101",  -- sqrt( 429) = 21
"000010101",  -- sqrt( 430) = 21
"000010101",  -- sqrt( 431) = 21
"000010101",  -- sqrt( 432) = 21
"000010101",  -- sqrt( 433) = 21
"000010101",  -- sqrt( 434) = 21
"000010101",  -- sqrt( 435) = 21
"000010101",  -- sqrt( 436) = 21
"000010101",  -- sqrt( 437) = 21
"000010101",  -- sqrt( 438) = 21
"000010101",  -- sqrt( 439) = 21
"000010101",  -- sqrt( 440) = 21
"000010101",  -- sqrt( 441) = 21
"000010101",  -- sqrt( 442) = 21
"000010101",  -- sqrt( 443) = 21
"000010101",  -- sqrt( 444) = 21
"000010101",  -- sqrt( 445) = 21
"000010101",  -- sqrt( 446) = 21
"000010101",  -- sqrt( 447) = 21
"000010101",  -- sqrt( 448) = 21
"000010101",  -- sqrt( 449) = 21
"000010101",  -- sqrt( 450) = 21
"000010101",  -- sqrt( 451) = 21
"000010101",  -- sqrt( 452) = 21
"000010101",  -- sqrt( 453) = 21
"000010101",  -- sqrt( 454) = 21
"000010101",  -- sqrt( 455) = 21
"000010101",  -- sqrt( 456) = 21
"000010101",  -- sqrt( 457) = 21
"000010101",  -- sqrt( 458) = 21
"000010101",  -- sqrt( 459) = 21
"000010101",  -- sqrt( 460) = 21
"000010101",  -- sqrt( 461) = 21
"000010101",  -- sqrt( 462) = 21
"000010110",  -- sqrt( 463) = 22
"000010110",  -- sqrt( 464) = 22
"000010110",  -- sqrt( 465) = 22
"000010110",  -- sqrt( 466) = 22
"000010110",  -- sqrt( 467) = 22
"000010110",  -- sqrt( 468) = 22
"000010110",  -- sqrt( 469) = 22
"000010110",  -- sqrt( 470) = 22
"000010110",  -- sqrt( 471) = 22
"000010110",  -- sqrt( 472) = 22
"000010110",  -- sqrt( 473) = 22
"000010110",  -- sqrt( 474) = 22
"000010110",  -- sqrt( 475) = 22
"000010110",  -- sqrt( 476) = 22
"000010110",  -- sqrt( 477) = 22
"000010110",  -- sqrt( 478) = 22
"000010110",  -- sqrt( 479) = 22
"000010110",  -- sqrt( 480) = 22
"000010110",  -- sqrt( 481) = 22
"000010110",  -- sqrt( 482) = 22
"000010110",  -- sqrt( 483) = 22
"000010110",  -- sqrt( 484) = 22
"000010110",  -- sqrt( 485) = 22
"000010110",  -- sqrt( 486) = 22
"000010110",  -- sqrt( 487) = 22
"000010110",  -- sqrt( 488) = 22
"000010110",  -- sqrt( 489) = 22
"000010110",  -- sqrt( 490) = 22
"000010110",  -- sqrt( 491) = 22
"000010110",  -- sqrt( 492) = 22
"000010110",  -- sqrt( 493) = 22
"000010110",  -- sqrt( 494) = 22
"000010110",  -- sqrt( 495) = 22
"000010110",  -- sqrt( 496) = 22
"000010110",  -- sqrt( 497) = 22
"000010110",  -- sqrt( 498) = 22
"000010110",  -- sqrt( 499) = 22
"000010110",  -- sqrt( 500) = 22
"000010110",  -- sqrt( 501) = 22
"000010110",  -- sqrt( 502) = 22
"000010110",  -- sqrt( 503) = 22
"000010110",  -- sqrt( 504) = 22
"000010110",  -- sqrt( 505) = 22
"000010110",  -- sqrt( 506) = 22
"000010111",  -- sqrt( 507) = 23
"000010111",  -- sqrt( 508) = 23
"000010111",  -- sqrt( 509) = 23
"000010111",  -- sqrt( 510) = 23
"000010111",  -- sqrt( 511) = 23
"000010111",  -- sqrt( 512) = 23
"000010111",  -- sqrt( 513) = 23
"000010111",  -- sqrt( 514) = 23
"000010111",  -- sqrt( 515) = 23
"000010111",  -- sqrt( 516) = 23
"000010111",  -- sqrt( 517) = 23
"000010111",  -- sqrt( 518) = 23
"000010111",  -- sqrt( 519) = 23
"000010111",  -- sqrt( 520) = 23
"000010111",  -- sqrt( 521) = 23
"000010111",  -- sqrt( 522) = 23
"000010111",  -- sqrt( 523) = 23
"000010111",  -- sqrt( 524) = 23
"000010111",  -- sqrt( 525) = 23
"000010111",  -- sqrt( 526) = 23
"000010111",  -- sqrt( 527) = 23
"000010111",  -- sqrt( 528) = 23
"000010111",  -- sqrt( 529) = 23
"000010111",  -- sqrt( 530) = 23
"000010111",  -- sqrt( 531) = 23
"000010111",  -- sqrt( 532) = 23
"000010111",  -- sqrt( 533) = 23
"000010111",  -- sqrt( 534) = 23
"000010111",  -- sqrt( 535) = 23
"000010111",  -- sqrt( 536) = 23
"000010111",  -- sqrt( 537) = 23
"000010111",  -- sqrt( 538) = 23
"000010111",  -- sqrt( 539) = 23
"000010111",  -- sqrt( 540) = 23
"000010111",  -- sqrt( 541) = 23
"000010111",  -- sqrt( 542) = 23
"000010111",  -- sqrt( 543) = 23
"000010111",  -- sqrt( 544) = 23
"000010111",  -- sqrt( 545) = 23
"000010111",  -- sqrt( 546) = 23
"000010111",  -- sqrt( 547) = 23
"000010111",  -- sqrt( 548) = 23
"000010111",  -- sqrt( 549) = 23
"000010111",  -- sqrt( 550) = 23
"000010111",  -- sqrt( 551) = 23
"000010111",  -- sqrt( 552) = 23
"000011000",  -- sqrt( 553) = 24
"000011000",  -- sqrt( 554) = 24
"000011000",  -- sqrt( 555) = 24
"000011000",  -- sqrt( 556) = 24
"000011000",  -- sqrt( 557) = 24
"000011000",  -- sqrt( 558) = 24
"000011000",  -- sqrt( 559) = 24
"000011000",  -- sqrt( 560) = 24
"000011000",  -- sqrt( 561) = 24
"000011000",  -- sqrt( 562) = 24
"000011000",  -- sqrt( 563) = 24
"000011000",  -- sqrt( 564) = 24
"000011000",  -- sqrt( 565) = 24
"000011000",  -- sqrt( 566) = 24
"000011000",  -- sqrt( 567) = 24
"000011000",  -- sqrt( 568) = 24
"000011000",  -- sqrt( 569) = 24
"000011000",  -- sqrt( 570) = 24
"000011000",  -- sqrt( 571) = 24
"000011000",  -- sqrt( 572) = 24
"000011000",  -- sqrt( 573) = 24
"000011000",  -- sqrt( 574) = 24
"000011000",  -- sqrt( 575) = 24
"000011000",  -- sqrt( 576) = 24
"000011000",  -- sqrt( 577) = 24
"000011000",  -- sqrt( 578) = 24
"000011000",  -- sqrt( 579) = 24
"000011000",  -- sqrt( 580) = 24
"000011000",  -- sqrt( 581) = 24
"000011000",  -- sqrt( 582) = 24
"000011000",  -- sqrt( 583) = 24
"000011000",  -- sqrt( 584) = 24
"000011000",  -- sqrt( 585) = 24
"000011000",  -- sqrt( 586) = 24
"000011000",  -- sqrt( 587) = 24
"000011000",  -- sqrt( 588) = 24
"000011000",  -- sqrt( 589) = 24
"000011000",  -- sqrt( 590) = 24
"000011000",  -- sqrt( 591) = 24
"000011000",  -- sqrt( 592) = 24
"000011000",  -- sqrt( 593) = 24
"000011000",  -- sqrt( 594) = 24
"000011000",  -- sqrt( 595) = 24
"000011000",  -- sqrt( 596) = 24
"000011000",  -- sqrt( 597) = 24
"000011000",  -- sqrt( 598) = 24
"000011000",  -- sqrt( 599) = 24
"000011000",  -- sqrt( 600) = 24
"000011001",  -- sqrt( 601) = 25
"000011001",  -- sqrt( 602) = 25
"000011001",  -- sqrt( 603) = 25
"000011001",  -- sqrt( 604) = 25
"000011001",  -- sqrt( 605) = 25
"000011001",  -- sqrt( 606) = 25
"000011001",  -- sqrt( 607) = 25
"000011001",  -- sqrt( 608) = 25
"000011001",  -- sqrt( 609) = 25
"000011001",  -- sqrt( 610) = 25
"000011001",  -- sqrt( 611) = 25
"000011001",  -- sqrt( 612) = 25
"000011001",  -- sqrt( 613) = 25
"000011001",  -- sqrt( 614) = 25
"000011001",  -- sqrt( 615) = 25
"000011001",  -- sqrt( 616) = 25
"000011001",  -- sqrt( 617) = 25
"000011001",  -- sqrt( 618) = 25
"000011001",  -- sqrt( 619) = 25
"000011001",  -- sqrt( 620) = 25
"000011001",  -- sqrt( 621) = 25
"000011001",  -- sqrt( 622) = 25
"000011001",  -- sqrt( 623) = 25
"000011001",  -- sqrt( 624) = 25
"000011001",  -- sqrt( 625) = 25
"000011001",  -- sqrt( 626) = 25
"000011001",  -- sqrt( 627) = 25
"000011001",  -- sqrt( 628) = 25
"000011001",  -- sqrt( 629) = 25
"000011001",  -- sqrt( 630) = 25
"000011001",  -- sqrt( 631) = 25
"000011001",  -- sqrt( 632) = 25
"000011001",  -- sqrt( 633) = 25
"000011001",  -- sqrt( 634) = 25
"000011001",  -- sqrt( 635) = 25
"000011001",  -- sqrt( 636) = 25
"000011001",  -- sqrt( 637) = 25
"000011001",  -- sqrt( 638) = 25
"000011001",  -- sqrt( 639) = 25
"000011001",  -- sqrt( 640) = 25
"000011001",  -- sqrt( 641) = 25
"000011001",  -- sqrt( 642) = 25
"000011001",  -- sqrt( 643) = 25
"000011001",  -- sqrt( 644) = 25
"000011001",  -- sqrt( 645) = 25
"000011001",  -- sqrt( 646) = 25
"000011001",  -- sqrt( 647) = 25
"000011001",  -- sqrt( 648) = 25
"000011001",  -- sqrt( 649) = 25
"000011001",  -- sqrt( 650) = 25
"000011010",  -- sqrt( 651) = 26
"000011010",  -- sqrt( 652) = 26
"000011010",  -- sqrt( 653) = 26
"000011010",  -- sqrt( 654) = 26
"000011010",  -- sqrt( 655) = 26
"000011010",  -- sqrt( 656) = 26
"000011010",  -- sqrt( 657) = 26
"000011010",  -- sqrt( 658) = 26
"000011010",  -- sqrt( 659) = 26
"000011010",  -- sqrt( 660) = 26
"000011010",  -- sqrt( 661) = 26
"000011010",  -- sqrt( 662) = 26
"000011010",  -- sqrt( 663) = 26
"000011010",  -- sqrt( 664) = 26
"000011010",  -- sqrt( 665) = 26
"000011010",  -- sqrt( 666) = 26
"000011010",  -- sqrt( 667) = 26
"000011010",  -- sqrt( 668) = 26
"000011010",  -- sqrt( 669) = 26
"000011010",  -- sqrt( 670) = 26
"000011010",  -- sqrt( 671) = 26
"000011010",  -- sqrt( 672) = 26
"000011010",  -- sqrt( 673) = 26
"000011010",  -- sqrt( 674) = 26
"000011010",  -- sqrt( 675) = 26
"000011010",  -- sqrt( 676) = 26
"000011010",  -- sqrt( 677) = 26
"000011010",  -- sqrt( 678) = 26
"000011010",  -- sqrt( 679) = 26
"000011010",  -- sqrt( 680) = 26
"000011010",  -- sqrt( 681) = 26
"000011010",  -- sqrt( 682) = 26
"000011010",  -- sqrt( 683) = 26
"000011010",  -- sqrt( 684) = 26
"000011010",  -- sqrt( 685) = 26
"000011010",  -- sqrt( 686) = 26
"000011010",  -- sqrt( 687) = 26
"000011010",  -- sqrt( 688) = 26
"000011010",  -- sqrt( 689) = 26
"000011010",  -- sqrt( 690) = 26
"000011010",  -- sqrt( 691) = 26
"000011010",  -- sqrt( 692) = 26
"000011010",  -- sqrt( 693) = 26
"000011010",  -- sqrt( 694) = 26
"000011010",  -- sqrt( 695) = 26
"000011010",  -- sqrt( 696) = 26
"000011010",  -- sqrt( 697) = 26
"000011010",  -- sqrt( 698) = 26
"000011010",  -- sqrt( 699) = 26
"000011010",  -- sqrt( 700) = 26
"000011010",  -- sqrt( 701) = 26
"000011010",  -- sqrt( 702) = 26
"000011011",  -- sqrt( 703) = 27
"000011011",  -- sqrt( 704) = 27
"000011011",  -- sqrt( 705) = 27
"000011011",  -- sqrt( 706) = 27
"000011011",  -- sqrt( 707) = 27
"000011011",  -- sqrt( 708) = 27
"000011011",  -- sqrt( 709) = 27
"000011011",  -- sqrt( 710) = 27
"000011011",  -- sqrt( 711) = 27
"000011011",  -- sqrt( 712) = 27
"000011011",  -- sqrt( 713) = 27
"000011011",  -- sqrt( 714) = 27
"000011011",  -- sqrt( 715) = 27
"000011011",  -- sqrt( 716) = 27
"000011011",  -- sqrt( 717) = 27
"000011011",  -- sqrt( 718) = 27
"000011011",  -- sqrt( 719) = 27
"000011011",  -- sqrt( 720) = 27
"000011011",  -- sqrt( 721) = 27
"000011011",  -- sqrt( 722) = 27
"000011011",  -- sqrt( 723) = 27
"000011011",  -- sqrt( 724) = 27
"000011011",  -- sqrt( 725) = 27
"000011011",  -- sqrt( 726) = 27
"000011011",  -- sqrt( 727) = 27
"000011011",  -- sqrt( 728) = 27
"000011011",  -- sqrt( 729) = 27
"000011011",  -- sqrt( 730) = 27
"000011011",  -- sqrt( 731) = 27
"000011011",  -- sqrt( 732) = 27
"000011011",  -- sqrt( 733) = 27
"000011011",  -- sqrt( 734) = 27
"000011011",  -- sqrt( 735) = 27
"000011011",  -- sqrt( 736) = 27
"000011011",  -- sqrt( 737) = 27
"000011011",  -- sqrt( 738) = 27
"000011011",  -- sqrt( 739) = 27
"000011011",  -- sqrt( 740) = 27
"000011011",  -- sqrt( 741) = 27
"000011011",  -- sqrt( 742) = 27
"000011011",  -- sqrt( 743) = 27
"000011011",  -- sqrt( 744) = 27
"000011011",  -- sqrt( 745) = 27
"000011011",  -- sqrt( 746) = 27
"000011011",  -- sqrt( 747) = 27
"000011011",  -- sqrt( 748) = 27
"000011011",  -- sqrt( 749) = 27
"000011011",  -- sqrt( 750) = 27
"000011011",  -- sqrt( 751) = 27
"000011011",  -- sqrt( 752) = 27
"000011011",  -- sqrt( 753) = 27
"000011011",  -- sqrt( 754) = 27
"000011011",  -- sqrt( 755) = 27
"000011011",  -- sqrt( 756) = 27
"000011100",  -- sqrt( 757) = 28
"000011100",  -- sqrt( 758) = 28
"000011100",  -- sqrt( 759) = 28
"000011100",  -- sqrt( 760) = 28
"000011100",  -- sqrt( 761) = 28
"000011100",  -- sqrt( 762) = 28
"000011100",  -- sqrt( 763) = 28
"000011100",  -- sqrt( 764) = 28
"000011100",  -- sqrt( 765) = 28
"000011100",  -- sqrt( 766) = 28
"000011100",  -- sqrt( 767) = 28
"000011100",  -- sqrt( 768) = 28
"000011100",  -- sqrt( 769) = 28
"000011100",  -- sqrt( 770) = 28
"000011100",  -- sqrt( 771) = 28
"000011100",  -- sqrt( 772) = 28
"000011100",  -- sqrt( 773) = 28
"000011100",  -- sqrt( 774) = 28
"000011100",  -- sqrt( 775) = 28
"000011100",  -- sqrt( 776) = 28
"000011100",  -- sqrt( 777) = 28
"000011100",  -- sqrt( 778) = 28
"000011100",  -- sqrt( 779) = 28
"000011100",  -- sqrt( 780) = 28
"000011100",  -- sqrt( 781) = 28
"000011100",  -- sqrt( 782) = 28
"000011100",  -- sqrt( 783) = 28
"000011100",  -- sqrt( 784) = 28
"000011100",  -- sqrt( 785) = 28
"000011100",  -- sqrt( 786) = 28
"000011100",  -- sqrt( 787) = 28
"000011100",  -- sqrt( 788) = 28
"000011100",  -- sqrt( 789) = 28
"000011100",  -- sqrt( 790) = 28
"000011100",  -- sqrt( 791) = 28
"000011100",  -- sqrt( 792) = 28
"000011100",  -- sqrt( 793) = 28
"000011100",  -- sqrt( 794) = 28
"000011100",  -- sqrt( 795) = 28
"000011100",  -- sqrt( 796) = 28
"000011100",  -- sqrt( 797) = 28
"000011100",  -- sqrt( 798) = 28
"000011100",  -- sqrt( 799) = 28
"000011100",  -- sqrt( 800) = 28
"000011100",  -- sqrt( 801) = 28
"000011100",  -- sqrt( 802) = 28
"000011100",  -- sqrt( 803) = 28
"000011100",  -- sqrt( 804) = 28
"000011100",  -- sqrt( 805) = 28
"000011100",  -- sqrt( 806) = 28
"000011100",  -- sqrt( 807) = 28
"000011100",  -- sqrt( 808) = 28
"000011100",  -- sqrt( 809) = 28
"000011100",  -- sqrt( 810) = 28
"000011100",  -- sqrt( 811) = 28
"000011100",  -- sqrt( 812) = 28
"000011101",  -- sqrt( 813) = 29
"000011101",  -- sqrt( 814) = 29
"000011101",  -- sqrt( 815) = 29
"000011101",  -- sqrt( 816) = 29
"000011101",  -- sqrt( 817) = 29
"000011101",  -- sqrt( 818) = 29
"000011101",  -- sqrt( 819) = 29
"000011101",  -- sqrt( 820) = 29
"000011101",  -- sqrt( 821) = 29
"000011101",  -- sqrt( 822) = 29
"000011101",  -- sqrt( 823) = 29
"000011101",  -- sqrt( 824) = 29
"000011101",  -- sqrt( 825) = 29
"000011101",  -- sqrt( 826) = 29
"000011101",  -- sqrt( 827) = 29
"000011101",  -- sqrt( 828) = 29
"000011101",  -- sqrt( 829) = 29
"000011101",  -- sqrt( 830) = 29
"000011101",  -- sqrt( 831) = 29
"000011101",  -- sqrt( 832) = 29
"000011101",  -- sqrt( 833) = 29
"000011101",  -- sqrt( 834) = 29
"000011101",  -- sqrt( 835) = 29
"000011101",  -- sqrt( 836) = 29
"000011101",  -- sqrt( 837) = 29
"000011101",  -- sqrt( 838) = 29
"000011101",  -- sqrt( 839) = 29
"000011101",  -- sqrt( 840) = 29
"000011101",  -- sqrt( 841) = 29
"000011101",  -- sqrt( 842) = 29
"000011101",  -- sqrt( 843) = 29
"000011101",  -- sqrt( 844) = 29
"000011101",  -- sqrt( 845) = 29
"000011101",  -- sqrt( 846) = 29
"000011101",  -- sqrt( 847) = 29
"000011101",  -- sqrt( 848) = 29
"000011101",  -- sqrt( 849) = 29
"000011101",  -- sqrt( 850) = 29
"000011101",  -- sqrt( 851) = 29
"000011101",  -- sqrt( 852) = 29
"000011101",  -- sqrt( 853) = 29
"000011101",  -- sqrt( 854) = 29
"000011101",  -- sqrt( 855) = 29
"000011101",  -- sqrt( 856) = 29
"000011101",  -- sqrt( 857) = 29
"000011101",  -- sqrt( 858) = 29
"000011101",  -- sqrt( 859) = 29
"000011101",  -- sqrt( 860) = 29
"000011101",  -- sqrt( 861) = 29
"000011101",  -- sqrt( 862) = 29
"000011101",  -- sqrt( 863) = 29
"000011101",  -- sqrt( 864) = 29
"000011101",  -- sqrt( 865) = 29
"000011101",  -- sqrt( 866) = 29
"000011101",  -- sqrt( 867) = 29
"000011101",  -- sqrt( 868) = 29
"000011101",  -- sqrt( 869) = 29
"000011101",  -- sqrt( 870) = 29
"000011110",  -- sqrt( 871) = 30
"000011110",  -- sqrt( 872) = 30
"000011110",  -- sqrt( 873) = 30
"000011110",  -- sqrt( 874) = 30
"000011110",  -- sqrt( 875) = 30
"000011110",  -- sqrt( 876) = 30
"000011110",  -- sqrt( 877) = 30
"000011110",  -- sqrt( 878) = 30
"000011110",  -- sqrt( 879) = 30
"000011110",  -- sqrt( 880) = 30
"000011110",  -- sqrt( 881) = 30
"000011110",  -- sqrt( 882) = 30
"000011110",  -- sqrt( 883) = 30
"000011110",  -- sqrt( 884) = 30
"000011110",  -- sqrt( 885) = 30
"000011110",  -- sqrt( 886) = 30
"000011110",  -- sqrt( 887) = 30
"000011110",  -- sqrt( 888) = 30
"000011110",  -- sqrt( 889) = 30
"000011110",  -- sqrt( 890) = 30
"000011110",  -- sqrt( 891) = 30
"000011110",  -- sqrt( 892) = 30
"000011110",  -- sqrt( 893) = 30
"000011110",  -- sqrt( 894) = 30
"000011110",  -- sqrt( 895) = 30
"000011110",  -- sqrt( 896) = 30
"000011110",  -- sqrt( 897) = 30
"000011110",  -- sqrt( 898) = 30
"000011110",  -- sqrt( 899) = 30
"000011110",  -- sqrt( 900) = 30
"000011110",  -- sqrt( 901) = 30
"000011110",  -- sqrt( 902) = 30
"000011110",  -- sqrt( 903) = 30
"000011110",  -- sqrt( 904) = 30
"000011110",  -- sqrt( 905) = 30
"000011110",  -- sqrt( 906) = 30
"000011110",  -- sqrt( 907) = 30
"000011110",  -- sqrt( 908) = 30
"000011110",  -- sqrt( 909) = 30
"000011110",  -- sqrt( 910) = 30
"000011110",  -- sqrt( 911) = 30
"000011110",  -- sqrt( 912) = 30
"000011110",  -- sqrt( 913) = 30
"000011110",  -- sqrt( 914) = 30
"000011110",  -- sqrt( 915) = 30
"000011110",  -- sqrt( 916) = 30
"000011110",  -- sqrt( 917) = 30
"000011110",  -- sqrt( 918) = 30
"000011110",  -- sqrt( 919) = 30
"000011110",  -- sqrt( 920) = 30
"000011110",  -- sqrt( 921) = 30
"000011110",  -- sqrt( 922) = 30
"000011110",  -- sqrt( 923) = 30
"000011110",  -- sqrt( 924) = 30
"000011110",  -- sqrt( 925) = 30
"000011110",  -- sqrt( 926) = 30
"000011110",  -- sqrt( 927) = 30
"000011110",  -- sqrt( 928) = 30
"000011110",  -- sqrt( 929) = 30
"000011110",  -- sqrt( 930) = 30
"000011111",  -- sqrt( 931) = 31
"000011111",  -- sqrt( 932) = 31
"000011111",  -- sqrt( 933) = 31
"000011111",  -- sqrt( 934) = 31
"000011111",  -- sqrt( 935) = 31
"000011111",  -- sqrt( 936) = 31
"000011111",  -- sqrt( 937) = 31
"000011111",  -- sqrt( 938) = 31
"000011111",  -- sqrt( 939) = 31
"000011111",  -- sqrt( 940) = 31
"000011111",  -- sqrt( 941) = 31
"000011111",  -- sqrt( 942) = 31
"000011111",  -- sqrt( 943) = 31
"000011111",  -- sqrt( 944) = 31
"000011111",  -- sqrt( 945) = 31
"000011111",  -- sqrt( 946) = 31
"000011111",  -- sqrt( 947) = 31
"000011111",  -- sqrt( 948) = 31
"000011111",  -- sqrt( 949) = 31
"000011111",  -- sqrt( 950) = 31
"000011111",  -- sqrt( 951) = 31
"000011111",  -- sqrt( 952) = 31
"000011111",  -- sqrt( 953) = 31
"000011111",  -- sqrt( 954) = 31
"000011111",  -- sqrt( 955) = 31
"000011111",  -- sqrt( 956) = 31
"000011111",  -- sqrt( 957) = 31
"000011111",  -- sqrt( 958) = 31
"000011111",  -- sqrt( 959) = 31
"000011111",  -- sqrt( 960) = 31
"000011111",  -- sqrt( 961) = 31
"000011111",  -- sqrt( 962) = 31
"000011111",  -- sqrt( 963) = 31
"000011111",  -- sqrt( 964) = 31
"000011111",  -- sqrt( 965) = 31
"000011111",  -- sqrt( 966) = 31
"000011111",  -- sqrt( 967) = 31
"000011111",  -- sqrt( 968) = 31
"000011111",  -- sqrt( 969) = 31
"000011111",  -- sqrt( 970) = 31
"000011111",  -- sqrt( 971) = 31
"000011111",  -- sqrt( 972) = 31
"000011111",  -- sqrt( 973) = 31
"000011111",  -- sqrt( 974) = 31
"000011111",  -- sqrt( 975) = 31
"000011111",  -- sqrt( 976) = 31
"000011111",  -- sqrt( 977) = 31
"000011111",  -- sqrt( 978) = 31
"000011111",  -- sqrt( 979) = 31
"000011111",  -- sqrt( 980) = 31
"000011111",  -- sqrt( 981) = 31
"000011111",  -- sqrt( 982) = 31
"000011111",  -- sqrt( 983) = 31
"000011111",  -- sqrt( 984) = 31
"000011111",  -- sqrt( 985) = 31
"000011111",  -- sqrt( 986) = 31
"000011111",  -- sqrt( 987) = 31
"000011111",  -- sqrt( 988) = 31
"000011111",  -- sqrt( 989) = 31
"000011111",  -- sqrt( 990) = 31
"000011111",  -- sqrt( 991) = 31
"000011111",  -- sqrt( 992) = 31
"000100000",  -- sqrt( 993) = 32
"000100000",  -- sqrt( 994) = 32
"000100000",  -- sqrt( 995) = 32
"000100000",  -- sqrt( 996) = 32
"000100000",  -- sqrt( 997) = 32
"000100000",  -- sqrt( 998) = 32
"000100000",  -- sqrt( 999) = 32
"000100000",  -- sqrt(1000) = 32
"000100000",  -- sqrt(1001) = 32
"000100000",  -- sqrt(1002) = 32
"000100000",  -- sqrt(1003) = 32
"000100000",  -- sqrt(1004) = 32
"000100000",  -- sqrt(1005) = 32
"000100000",  -- sqrt(1006) = 32
"000100000",  -- sqrt(1007) = 32
"000100000",  -- sqrt(1008) = 32
"000100000",  -- sqrt(1009) = 32
"000100000",  -- sqrt(1010) = 32
"000100000",  -- sqrt(1011) = 32
"000100000",  -- sqrt(1012) = 32
"000100000",  -- sqrt(1013) = 32
"000100000",  -- sqrt(1014) = 32
"000100000",  -- sqrt(1015) = 32
"000100000",  -- sqrt(1016) = 32
"000100000",  -- sqrt(1017) = 32
"000100000",  -- sqrt(1018) = 32
"000100000",  -- sqrt(1019) = 32
"000100000",  -- sqrt(1020) = 32
"000100000",  -- sqrt(1021) = 32
"000100000",  -- sqrt(1022) = 32
"000100000",  -- sqrt(1023) = 32
"000100000",  -- sqrt(1024) = 32
"000100000",  -- sqrt(1025) = 32
"000100000",  -- sqrt(1026) = 32
"000100000",  -- sqrt(1027) = 32
"000100000",  -- sqrt(1028) = 32
"000100000",  -- sqrt(1029) = 32
"000100000",  -- sqrt(1030) = 32
"000100000",  -- sqrt(1031) = 32
"000100000",  -- sqrt(1032) = 32
"000100000",  -- sqrt(1033) = 32
"000100000",  -- sqrt(1034) = 32
"000100000",  -- sqrt(1035) = 32
"000100000",  -- sqrt(1036) = 32
"000100000",  -- sqrt(1037) = 32
"000100000",  -- sqrt(1038) = 32
"000100000",  -- sqrt(1039) = 32
"000100000",  -- sqrt(1040) = 32
"000100000",  -- sqrt(1041) = 32
"000100000",  -- sqrt(1042) = 32
"000100000",  -- sqrt(1043) = 32
"000100000",  -- sqrt(1044) = 32
"000100000",  -- sqrt(1045) = 32
"000100000",  -- sqrt(1046) = 32
"000100000",  -- sqrt(1047) = 32
"000100000",  -- sqrt(1048) = 32
"000100000",  -- sqrt(1049) = 32
"000100000",  -- sqrt(1050) = 32
"000100000",  -- sqrt(1051) = 32
"000100000",  -- sqrt(1052) = 32
"000100000",  -- sqrt(1053) = 32
"000100000",  -- sqrt(1054) = 32
"000100000",  -- sqrt(1055) = 32
"000100000",  -- sqrt(1056) = 32
"000100001",  -- sqrt(1057) = 33
"000100001",  -- sqrt(1058) = 33
"000100001",  -- sqrt(1059) = 33
"000100001",  -- sqrt(1060) = 33
"000100001",  -- sqrt(1061) = 33
"000100001",  -- sqrt(1062) = 33
"000100001",  -- sqrt(1063) = 33
"000100001",  -- sqrt(1064) = 33
"000100001",  -- sqrt(1065) = 33
"000100001",  -- sqrt(1066) = 33
"000100001",  -- sqrt(1067) = 33
"000100001",  -- sqrt(1068) = 33
"000100001",  -- sqrt(1069) = 33
"000100001",  -- sqrt(1070) = 33
"000100001",  -- sqrt(1071) = 33
"000100001",  -- sqrt(1072) = 33
"000100001",  -- sqrt(1073) = 33
"000100001",  -- sqrt(1074) = 33
"000100001",  -- sqrt(1075) = 33
"000100001",  -- sqrt(1076) = 33
"000100001",  -- sqrt(1077) = 33
"000100001",  -- sqrt(1078) = 33
"000100001",  -- sqrt(1079) = 33
"000100001",  -- sqrt(1080) = 33
"000100001",  -- sqrt(1081) = 33
"000100001",  -- sqrt(1082) = 33
"000100001",  -- sqrt(1083) = 33
"000100001",  -- sqrt(1084) = 33
"000100001",  -- sqrt(1085) = 33
"000100001",  -- sqrt(1086) = 33
"000100001",  -- sqrt(1087) = 33
"000100001",  -- sqrt(1088) = 33
"000100001",  -- sqrt(1089) = 33
"000100001",  -- sqrt(1090) = 33
"000100001",  -- sqrt(1091) = 33
"000100001",  -- sqrt(1092) = 33
"000100001",  -- sqrt(1093) = 33
"000100001",  -- sqrt(1094) = 33
"000100001",  -- sqrt(1095) = 33
"000100001",  -- sqrt(1096) = 33
"000100001",  -- sqrt(1097) = 33
"000100001",  -- sqrt(1098) = 33
"000100001",  -- sqrt(1099) = 33
"000100001",  -- sqrt(1100) = 33
"000100001",  -- sqrt(1101) = 33
"000100001",  -- sqrt(1102) = 33
"000100001",  -- sqrt(1103) = 33
"000100001",  -- sqrt(1104) = 33
"000100001",  -- sqrt(1105) = 33
"000100001",  -- sqrt(1106) = 33
"000100001",  -- sqrt(1107) = 33
"000100001",  -- sqrt(1108) = 33
"000100001",  -- sqrt(1109) = 33
"000100001",  -- sqrt(1110) = 33
"000100001",  -- sqrt(1111) = 33
"000100001",  -- sqrt(1112) = 33
"000100001",  -- sqrt(1113) = 33
"000100001",  -- sqrt(1114) = 33
"000100001",  -- sqrt(1115) = 33
"000100001",  -- sqrt(1116) = 33
"000100001",  -- sqrt(1117) = 33
"000100001",  -- sqrt(1118) = 33
"000100001",  -- sqrt(1119) = 33
"000100001",  -- sqrt(1120) = 33
"000100001",  -- sqrt(1121) = 33
"000100001",  -- sqrt(1122) = 33
"000100010",  -- sqrt(1123) = 34
"000100010",  -- sqrt(1124) = 34
"000100010",  -- sqrt(1125) = 34
"000100010",  -- sqrt(1126) = 34
"000100010",  -- sqrt(1127) = 34
"000100010",  -- sqrt(1128) = 34
"000100010",  -- sqrt(1129) = 34
"000100010",  -- sqrt(1130) = 34
"000100010",  -- sqrt(1131) = 34
"000100010",  -- sqrt(1132) = 34
"000100010",  -- sqrt(1133) = 34
"000100010",  -- sqrt(1134) = 34
"000100010",  -- sqrt(1135) = 34
"000100010",  -- sqrt(1136) = 34
"000100010",  -- sqrt(1137) = 34
"000100010",  -- sqrt(1138) = 34
"000100010",  -- sqrt(1139) = 34
"000100010",  -- sqrt(1140) = 34
"000100010",  -- sqrt(1141) = 34
"000100010",  -- sqrt(1142) = 34
"000100010",  -- sqrt(1143) = 34
"000100010",  -- sqrt(1144) = 34
"000100010",  -- sqrt(1145) = 34
"000100010",  -- sqrt(1146) = 34
"000100010",  -- sqrt(1147) = 34
"000100010",  -- sqrt(1148) = 34
"000100010",  -- sqrt(1149) = 34
"000100010",  -- sqrt(1150) = 34
"000100010",  -- sqrt(1151) = 34
"000100010",  -- sqrt(1152) = 34
"000100010",  -- sqrt(1153) = 34
"000100010",  -- sqrt(1154) = 34
"000100010",  -- sqrt(1155) = 34
"000100010",  -- sqrt(1156) = 34
"000100010",  -- sqrt(1157) = 34
"000100010",  -- sqrt(1158) = 34
"000100010",  -- sqrt(1159) = 34
"000100010",  -- sqrt(1160) = 34
"000100010",  -- sqrt(1161) = 34
"000100010",  -- sqrt(1162) = 34
"000100010",  -- sqrt(1163) = 34
"000100010",  -- sqrt(1164) = 34
"000100010",  -- sqrt(1165) = 34
"000100010",  -- sqrt(1166) = 34
"000100010",  -- sqrt(1167) = 34
"000100010",  -- sqrt(1168) = 34
"000100010",  -- sqrt(1169) = 34
"000100010",  -- sqrt(1170) = 34
"000100010",  -- sqrt(1171) = 34
"000100010",  -- sqrt(1172) = 34
"000100010",  -- sqrt(1173) = 34
"000100010",  -- sqrt(1174) = 34
"000100010",  -- sqrt(1175) = 34
"000100010",  -- sqrt(1176) = 34
"000100010",  -- sqrt(1177) = 34
"000100010",  -- sqrt(1178) = 34
"000100010",  -- sqrt(1179) = 34
"000100010",  -- sqrt(1180) = 34
"000100010",  -- sqrt(1181) = 34
"000100010",  -- sqrt(1182) = 34
"000100010",  -- sqrt(1183) = 34
"000100010",  -- sqrt(1184) = 34
"000100010",  -- sqrt(1185) = 34
"000100010",  -- sqrt(1186) = 34
"000100010",  -- sqrt(1187) = 34
"000100010",  -- sqrt(1188) = 34
"000100010",  -- sqrt(1189) = 34
"000100010",  -- sqrt(1190) = 34
"000100011",  -- sqrt(1191) = 35
"000100011",  -- sqrt(1192) = 35
"000100011",  -- sqrt(1193) = 35
"000100011",  -- sqrt(1194) = 35
"000100011",  -- sqrt(1195) = 35
"000100011",  -- sqrt(1196) = 35
"000100011",  -- sqrt(1197) = 35
"000100011",  -- sqrt(1198) = 35
"000100011",  -- sqrt(1199) = 35
"000100011",  -- sqrt(1200) = 35
"000100011",  -- sqrt(1201) = 35
"000100011",  -- sqrt(1202) = 35
"000100011",  -- sqrt(1203) = 35
"000100011",  -- sqrt(1204) = 35
"000100011",  -- sqrt(1205) = 35
"000100011",  -- sqrt(1206) = 35
"000100011",  -- sqrt(1207) = 35
"000100011",  -- sqrt(1208) = 35
"000100011",  -- sqrt(1209) = 35
"000100011",  -- sqrt(1210) = 35
"000100011",  -- sqrt(1211) = 35
"000100011",  -- sqrt(1212) = 35
"000100011",  -- sqrt(1213) = 35
"000100011",  -- sqrt(1214) = 35
"000100011",  -- sqrt(1215) = 35
"000100011",  -- sqrt(1216) = 35
"000100011",  -- sqrt(1217) = 35
"000100011",  -- sqrt(1218) = 35
"000100011",  -- sqrt(1219) = 35
"000100011",  -- sqrt(1220) = 35
"000100011",  -- sqrt(1221) = 35
"000100011",  -- sqrt(1222) = 35
"000100011",  -- sqrt(1223) = 35
"000100011",  -- sqrt(1224) = 35
"000100011",  -- sqrt(1225) = 35
"000100011",  -- sqrt(1226) = 35
"000100011",  -- sqrt(1227) = 35
"000100011",  -- sqrt(1228) = 35
"000100011",  -- sqrt(1229) = 35
"000100011",  -- sqrt(1230) = 35
"000100011",  -- sqrt(1231) = 35
"000100011",  -- sqrt(1232) = 35
"000100011",  -- sqrt(1233) = 35
"000100011",  -- sqrt(1234) = 35
"000100011",  -- sqrt(1235) = 35
"000100011",  -- sqrt(1236) = 35
"000100011",  -- sqrt(1237) = 35
"000100011",  -- sqrt(1238) = 35
"000100011",  -- sqrt(1239) = 35
"000100011",  -- sqrt(1240) = 35
"000100011",  -- sqrt(1241) = 35
"000100011",  -- sqrt(1242) = 35
"000100011",  -- sqrt(1243) = 35
"000100011",  -- sqrt(1244) = 35
"000100011",  -- sqrt(1245) = 35
"000100011",  -- sqrt(1246) = 35
"000100011",  -- sqrt(1247) = 35
"000100011",  -- sqrt(1248) = 35
"000100011",  -- sqrt(1249) = 35
"000100011",  -- sqrt(1250) = 35
"000100011",  -- sqrt(1251) = 35
"000100011",  -- sqrt(1252) = 35
"000100011",  -- sqrt(1253) = 35
"000100011",  -- sqrt(1254) = 35
"000100011",  -- sqrt(1255) = 35
"000100011",  -- sqrt(1256) = 35
"000100011",  -- sqrt(1257) = 35
"000100011",  -- sqrt(1258) = 35
"000100011",  -- sqrt(1259) = 35
"000100011",  -- sqrt(1260) = 35
"000100100",  -- sqrt(1261) = 36
"000100100",  -- sqrt(1262) = 36
"000100100",  -- sqrt(1263) = 36
"000100100",  -- sqrt(1264) = 36
"000100100",  -- sqrt(1265) = 36
"000100100",  -- sqrt(1266) = 36
"000100100",  -- sqrt(1267) = 36
"000100100",  -- sqrt(1268) = 36
"000100100",  -- sqrt(1269) = 36
"000100100",  -- sqrt(1270) = 36
"000100100",  -- sqrt(1271) = 36
"000100100",  -- sqrt(1272) = 36
"000100100",  -- sqrt(1273) = 36
"000100100",  -- sqrt(1274) = 36
"000100100",  -- sqrt(1275) = 36
"000100100",  -- sqrt(1276) = 36
"000100100",  -- sqrt(1277) = 36
"000100100",  -- sqrt(1278) = 36
"000100100",  -- sqrt(1279) = 36
"000100100",  -- sqrt(1280) = 36
"000100100",  -- sqrt(1281) = 36
"000100100",  -- sqrt(1282) = 36
"000100100",  -- sqrt(1283) = 36
"000100100",  -- sqrt(1284) = 36
"000100100",  -- sqrt(1285) = 36
"000100100",  -- sqrt(1286) = 36
"000100100",  -- sqrt(1287) = 36
"000100100",  -- sqrt(1288) = 36
"000100100",  -- sqrt(1289) = 36
"000100100",  -- sqrt(1290) = 36
"000100100",  -- sqrt(1291) = 36
"000100100",  -- sqrt(1292) = 36
"000100100",  -- sqrt(1293) = 36
"000100100",  -- sqrt(1294) = 36
"000100100",  -- sqrt(1295) = 36
"000100100",  -- sqrt(1296) = 36
"000100100",  -- sqrt(1297) = 36
"000100100",  -- sqrt(1298) = 36
"000100100",  -- sqrt(1299) = 36
"000100100",  -- sqrt(1300) = 36
"000100100",  -- sqrt(1301) = 36
"000100100",  -- sqrt(1302) = 36
"000100100",  -- sqrt(1303) = 36
"000100100",  -- sqrt(1304) = 36
"000100100",  -- sqrt(1305) = 36
"000100100",  -- sqrt(1306) = 36
"000100100",  -- sqrt(1307) = 36
"000100100",  -- sqrt(1308) = 36
"000100100",  -- sqrt(1309) = 36
"000100100",  -- sqrt(1310) = 36
"000100100",  -- sqrt(1311) = 36
"000100100",  -- sqrt(1312) = 36
"000100100",  -- sqrt(1313) = 36
"000100100",  -- sqrt(1314) = 36
"000100100",  -- sqrt(1315) = 36
"000100100",  -- sqrt(1316) = 36
"000100100",  -- sqrt(1317) = 36
"000100100",  -- sqrt(1318) = 36
"000100100",  -- sqrt(1319) = 36
"000100100",  -- sqrt(1320) = 36
"000100100",  -- sqrt(1321) = 36
"000100100",  -- sqrt(1322) = 36
"000100100",  -- sqrt(1323) = 36
"000100100",  -- sqrt(1324) = 36
"000100100",  -- sqrt(1325) = 36
"000100100",  -- sqrt(1326) = 36
"000100100",  -- sqrt(1327) = 36
"000100100",  -- sqrt(1328) = 36
"000100100",  -- sqrt(1329) = 36
"000100100",  -- sqrt(1330) = 36
"000100100",  -- sqrt(1331) = 36
"000100100",  -- sqrt(1332) = 36
"000100101",  -- sqrt(1333) = 37
"000100101",  -- sqrt(1334) = 37
"000100101",  -- sqrt(1335) = 37
"000100101",  -- sqrt(1336) = 37
"000100101",  -- sqrt(1337) = 37
"000100101",  -- sqrt(1338) = 37
"000100101",  -- sqrt(1339) = 37
"000100101",  -- sqrt(1340) = 37
"000100101",  -- sqrt(1341) = 37
"000100101",  -- sqrt(1342) = 37
"000100101",  -- sqrt(1343) = 37
"000100101",  -- sqrt(1344) = 37
"000100101",  -- sqrt(1345) = 37
"000100101",  -- sqrt(1346) = 37
"000100101",  -- sqrt(1347) = 37
"000100101",  -- sqrt(1348) = 37
"000100101",  -- sqrt(1349) = 37
"000100101",  -- sqrt(1350) = 37
"000100101",  -- sqrt(1351) = 37
"000100101",  -- sqrt(1352) = 37
"000100101",  -- sqrt(1353) = 37
"000100101",  -- sqrt(1354) = 37
"000100101",  -- sqrt(1355) = 37
"000100101",  -- sqrt(1356) = 37
"000100101",  -- sqrt(1357) = 37
"000100101",  -- sqrt(1358) = 37
"000100101",  -- sqrt(1359) = 37
"000100101",  -- sqrt(1360) = 37
"000100101",  -- sqrt(1361) = 37
"000100101",  -- sqrt(1362) = 37
"000100101",  -- sqrt(1363) = 37
"000100101",  -- sqrt(1364) = 37
"000100101",  -- sqrt(1365) = 37
"000100101",  -- sqrt(1366) = 37
"000100101",  -- sqrt(1367) = 37
"000100101",  -- sqrt(1368) = 37
"000100101",  -- sqrt(1369) = 37
"000100101",  -- sqrt(1370) = 37
"000100101",  -- sqrt(1371) = 37
"000100101",  -- sqrt(1372) = 37
"000100101",  -- sqrt(1373) = 37
"000100101",  -- sqrt(1374) = 37
"000100101",  -- sqrt(1375) = 37
"000100101",  -- sqrt(1376) = 37
"000100101",  -- sqrt(1377) = 37
"000100101",  -- sqrt(1378) = 37
"000100101",  -- sqrt(1379) = 37
"000100101",  -- sqrt(1380) = 37
"000100101",  -- sqrt(1381) = 37
"000100101",  -- sqrt(1382) = 37
"000100101",  -- sqrt(1383) = 37
"000100101",  -- sqrt(1384) = 37
"000100101",  -- sqrt(1385) = 37
"000100101",  -- sqrt(1386) = 37
"000100101",  -- sqrt(1387) = 37
"000100101",  -- sqrt(1388) = 37
"000100101",  -- sqrt(1389) = 37
"000100101",  -- sqrt(1390) = 37
"000100101",  -- sqrt(1391) = 37
"000100101",  -- sqrt(1392) = 37
"000100101",  -- sqrt(1393) = 37
"000100101",  -- sqrt(1394) = 37
"000100101",  -- sqrt(1395) = 37
"000100101",  -- sqrt(1396) = 37
"000100101",  -- sqrt(1397) = 37
"000100101",  -- sqrt(1398) = 37
"000100101",  -- sqrt(1399) = 37
"000100101",  -- sqrt(1400) = 37
"000100101",  -- sqrt(1401) = 37
"000100101",  -- sqrt(1402) = 37
"000100101",  -- sqrt(1403) = 37
"000100101",  -- sqrt(1404) = 37
"000100101",  -- sqrt(1405) = 37
"000100101",  -- sqrt(1406) = 37
"000100110",  -- sqrt(1407) = 38
"000100110",  -- sqrt(1408) = 38
"000100110",  -- sqrt(1409) = 38
"000100110",  -- sqrt(1410) = 38
"000100110",  -- sqrt(1411) = 38
"000100110",  -- sqrt(1412) = 38
"000100110",  -- sqrt(1413) = 38
"000100110",  -- sqrt(1414) = 38
"000100110",  -- sqrt(1415) = 38
"000100110",  -- sqrt(1416) = 38
"000100110",  -- sqrt(1417) = 38
"000100110",  -- sqrt(1418) = 38
"000100110",  -- sqrt(1419) = 38
"000100110",  -- sqrt(1420) = 38
"000100110",  -- sqrt(1421) = 38
"000100110",  -- sqrt(1422) = 38
"000100110",  -- sqrt(1423) = 38
"000100110",  -- sqrt(1424) = 38
"000100110",  -- sqrt(1425) = 38
"000100110",  -- sqrt(1426) = 38
"000100110",  -- sqrt(1427) = 38
"000100110",  -- sqrt(1428) = 38
"000100110",  -- sqrt(1429) = 38
"000100110",  -- sqrt(1430) = 38
"000100110",  -- sqrt(1431) = 38
"000100110",  -- sqrt(1432) = 38
"000100110",  -- sqrt(1433) = 38
"000100110",  -- sqrt(1434) = 38
"000100110",  -- sqrt(1435) = 38
"000100110",  -- sqrt(1436) = 38
"000100110",  -- sqrt(1437) = 38
"000100110",  -- sqrt(1438) = 38
"000100110",  -- sqrt(1439) = 38
"000100110",  -- sqrt(1440) = 38
"000100110",  -- sqrt(1441) = 38
"000100110",  -- sqrt(1442) = 38
"000100110",  -- sqrt(1443) = 38
"000100110",  -- sqrt(1444) = 38
"000100110",  -- sqrt(1445) = 38
"000100110",  -- sqrt(1446) = 38
"000100110",  -- sqrt(1447) = 38
"000100110",  -- sqrt(1448) = 38
"000100110",  -- sqrt(1449) = 38
"000100110",  -- sqrt(1450) = 38
"000100110",  -- sqrt(1451) = 38
"000100110",  -- sqrt(1452) = 38
"000100110",  -- sqrt(1453) = 38
"000100110",  -- sqrt(1454) = 38
"000100110",  -- sqrt(1455) = 38
"000100110",  -- sqrt(1456) = 38
"000100110",  -- sqrt(1457) = 38
"000100110",  -- sqrt(1458) = 38
"000100110",  -- sqrt(1459) = 38
"000100110",  -- sqrt(1460) = 38
"000100110",  -- sqrt(1461) = 38
"000100110",  -- sqrt(1462) = 38
"000100110",  -- sqrt(1463) = 38
"000100110",  -- sqrt(1464) = 38
"000100110",  -- sqrt(1465) = 38
"000100110",  -- sqrt(1466) = 38
"000100110",  -- sqrt(1467) = 38
"000100110",  -- sqrt(1468) = 38
"000100110",  -- sqrt(1469) = 38
"000100110",  -- sqrt(1470) = 38
"000100110",  -- sqrt(1471) = 38
"000100110",  -- sqrt(1472) = 38
"000100110",  -- sqrt(1473) = 38
"000100110",  -- sqrt(1474) = 38
"000100110",  -- sqrt(1475) = 38
"000100110",  -- sqrt(1476) = 38
"000100110",  -- sqrt(1477) = 38
"000100110",  -- sqrt(1478) = 38
"000100110",  -- sqrt(1479) = 38
"000100110",  -- sqrt(1480) = 38
"000100110",  -- sqrt(1481) = 38
"000100110",  -- sqrt(1482) = 38
"000100111",  -- sqrt(1483) = 39
"000100111",  -- sqrt(1484) = 39
"000100111",  -- sqrt(1485) = 39
"000100111",  -- sqrt(1486) = 39
"000100111",  -- sqrt(1487) = 39
"000100111",  -- sqrt(1488) = 39
"000100111",  -- sqrt(1489) = 39
"000100111",  -- sqrt(1490) = 39
"000100111",  -- sqrt(1491) = 39
"000100111",  -- sqrt(1492) = 39
"000100111",  -- sqrt(1493) = 39
"000100111",  -- sqrt(1494) = 39
"000100111",  -- sqrt(1495) = 39
"000100111",  -- sqrt(1496) = 39
"000100111",  -- sqrt(1497) = 39
"000100111",  -- sqrt(1498) = 39
"000100111",  -- sqrt(1499) = 39
"000100111",  -- sqrt(1500) = 39
"000100111",  -- sqrt(1501) = 39
"000100111",  -- sqrt(1502) = 39
"000100111",  -- sqrt(1503) = 39
"000100111",  -- sqrt(1504) = 39
"000100111",  -- sqrt(1505) = 39
"000100111",  -- sqrt(1506) = 39
"000100111",  -- sqrt(1507) = 39
"000100111",  -- sqrt(1508) = 39
"000100111",  -- sqrt(1509) = 39
"000100111",  -- sqrt(1510) = 39
"000100111",  -- sqrt(1511) = 39
"000100111",  -- sqrt(1512) = 39
"000100111",  -- sqrt(1513) = 39
"000100111",  -- sqrt(1514) = 39
"000100111",  -- sqrt(1515) = 39
"000100111",  -- sqrt(1516) = 39
"000100111",  -- sqrt(1517) = 39
"000100111",  -- sqrt(1518) = 39
"000100111",  -- sqrt(1519) = 39
"000100111",  -- sqrt(1520) = 39
"000100111",  -- sqrt(1521) = 39
"000100111",  -- sqrt(1522) = 39
"000100111",  -- sqrt(1523) = 39
"000100111",  -- sqrt(1524) = 39
"000100111",  -- sqrt(1525) = 39
"000100111",  -- sqrt(1526) = 39
"000100111",  -- sqrt(1527) = 39
"000100111",  -- sqrt(1528) = 39
"000100111",  -- sqrt(1529) = 39
"000100111",  -- sqrt(1530) = 39
"000100111",  -- sqrt(1531) = 39
"000100111",  -- sqrt(1532) = 39
"000100111",  -- sqrt(1533) = 39
"000100111",  -- sqrt(1534) = 39
"000100111",  -- sqrt(1535) = 39
"000100111",  -- sqrt(1536) = 39
"000100111",  -- sqrt(1537) = 39
"000100111",  -- sqrt(1538) = 39
"000100111",  -- sqrt(1539) = 39
"000100111",  -- sqrt(1540) = 39
"000100111",  -- sqrt(1541) = 39
"000100111",  -- sqrt(1542) = 39
"000100111",  -- sqrt(1543) = 39
"000100111",  -- sqrt(1544) = 39
"000100111",  -- sqrt(1545) = 39
"000100111",  -- sqrt(1546) = 39
"000100111",  -- sqrt(1547) = 39
"000100111",  -- sqrt(1548) = 39
"000100111",  -- sqrt(1549) = 39
"000100111",  -- sqrt(1550) = 39
"000100111",  -- sqrt(1551) = 39
"000100111",  -- sqrt(1552) = 39
"000100111",  -- sqrt(1553) = 39
"000100111",  -- sqrt(1554) = 39
"000100111",  -- sqrt(1555) = 39
"000100111",  -- sqrt(1556) = 39
"000100111",  -- sqrt(1557) = 39
"000100111",  -- sqrt(1558) = 39
"000100111",  -- sqrt(1559) = 39
"000100111",  -- sqrt(1560) = 39
"000101000",  -- sqrt(1561) = 40
"000101000",  -- sqrt(1562) = 40
"000101000",  -- sqrt(1563) = 40
"000101000",  -- sqrt(1564) = 40
"000101000",  -- sqrt(1565) = 40
"000101000",  -- sqrt(1566) = 40
"000101000",  -- sqrt(1567) = 40
"000101000",  -- sqrt(1568) = 40
"000101000",  -- sqrt(1569) = 40
"000101000",  -- sqrt(1570) = 40
"000101000",  -- sqrt(1571) = 40
"000101000",  -- sqrt(1572) = 40
"000101000",  -- sqrt(1573) = 40
"000101000",  -- sqrt(1574) = 40
"000101000",  -- sqrt(1575) = 40
"000101000",  -- sqrt(1576) = 40
"000101000",  -- sqrt(1577) = 40
"000101000",  -- sqrt(1578) = 40
"000101000",  -- sqrt(1579) = 40
"000101000",  -- sqrt(1580) = 40
"000101000",  -- sqrt(1581) = 40
"000101000",  -- sqrt(1582) = 40
"000101000",  -- sqrt(1583) = 40
"000101000",  -- sqrt(1584) = 40
"000101000",  -- sqrt(1585) = 40
"000101000",  -- sqrt(1586) = 40
"000101000",  -- sqrt(1587) = 40
"000101000",  -- sqrt(1588) = 40
"000101000",  -- sqrt(1589) = 40
"000101000",  -- sqrt(1590) = 40
"000101000",  -- sqrt(1591) = 40
"000101000",  -- sqrt(1592) = 40
"000101000",  -- sqrt(1593) = 40
"000101000",  -- sqrt(1594) = 40
"000101000",  -- sqrt(1595) = 40
"000101000",  -- sqrt(1596) = 40
"000101000",  -- sqrt(1597) = 40
"000101000",  -- sqrt(1598) = 40
"000101000",  -- sqrt(1599) = 40
"000101000",  -- sqrt(1600) = 40
"000101000",  -- sqrt(1601) = 40
"000101000",  -- sqrt(1602) = 40
"000101000",  -- sqrt(1603) = 40
"000101000",  -- sqrt(1604) = 40
"000101000",  -- sqrt(1605) = 40
"000101000",  -- sqrt(1606) = 40
"000101000",  -- sqrt(1607) = 40
"000101000",  -- sqrt(1608) = 40
"000101000",  -- sqrt(1609) = 40
"000101000",  -- sqrt(1610) = 40
"000101000",  -- sqrt(1611) = 40
"000101000",  -- sqrt(1612) = 40
"000101000",  -- sqrt(1613) = 40
"000101000",  -- sqrt(1614) = 40
"000101000",  -- sqrt(1615) = 40
"000101000",  -- sqrt(1616) = 40
"000101000",  -- sqrt(1617) = 40
"000101000",  -- sqrt(1618) = 40
"000101000",  -- sqrt(1619) = 40
"000101000",  -- sqrt(1620) = 40
"000101000",  -- sqrt(1621) = 40
"000101000",  -- sqrt(1622) = 40
"000101000",  -- sqrt(1623) = 40
"000101000",  -- sqrt(1624) = 40
"000101000",  -- sqrt(1625) = 40
"000101000",  -- sqrt(1626) = 40
"000101000",  -- sqrt(1627) = 40
"000101000",  -- sqrt(1628) = 40
"000101000",  -- sqrt(1629) = 40
"000101000",  -- sqrt(1630) = 40
"000101000",  -- sqrt(1631) = 40
"000101000",  -- sqrt(1632) = 40
"000101000",  -- sqrt(1633) = 40
"000101000",  -- sqrt(1634) = 40
"000101000",  -- sqrt(1635) = 40
"000101000",  -- sqrt(1636) = 40
"000101000",  -- sqrt(1637) = 40
"000101000",  -- sqrt(1638) = 40
"000101000",  -- sqrt(1639) = 40
"000101000",  -- sqrt(1640) = 40
"000101001",  -- sqrt(1641) = 41
"000101001",  -- sqrt(1642) = 41
"000101001",  -- sqrt(1643) = 41
"000101001",  -- sqrt(1644) = 41
"000101001",  -- sqrt(1645) = 41
"000101001",  -- sqrt(1646) = 41
"000101001",  -- sqrt(1647) = 41
"000101001",  -- sqrt(1648) = 41
"000101001",  -- sqrt(1649) = 41
"000101001",  -- sqrt(1650) = 41
"000101001",  -- sqrt(1651) = 41
"000101001",  -- sqrt(1652) = 41
"000101001",  -- sqrt(1653) = 41
"000101001",  -- sqrt(1654) = 41
"000101001",  -- sqrt(1655) = 41
"000101001",  -- sqrt(1656) = 41
"000101001",  -- sqrt(1657) = 41
"000101001",  -- sqrt(1658) = 41
"000101001",  -- sqrt(1659) = 41
"000101001",  -- sqrt(1660) = 41
"000101001",  -- sqrt(1661) = 41
"000101001",  -- sqrt(1662) = 41
"000101001",  -- sqrt(1663) = 41
"000101001",  -- sqrt(1664) = 41
"000101001",  -- sqrt(1665) = 41
"000101001",  -- sqrt(1666) = 41
"000101001",  -- sqrt(1667) = 41
"000101001",  -- sqrt(1668) = 41
"000101001",  -- sqrt(1669) = 41
"000101001",  -- sqrt(1670) = 41
"000101001",  -- sqrt(1671) = 41
"000101001",  -- sqrt(1672) = 41
"000101001",  -- sqrt(1673) = 41
"000101001",  -- sqrt(1674) = 41
"000101001",  -- sqrt(1675) = 41
"000101001",  -- sqrt(1676) = 41
"000101001",  -- sqrt(1677) = 41
"000101001",  -- sqrt(1678) = 41
"000101001",  -- sqrt(1679) = 41
"000101001",  -- sqrt(1680) = 41
"000101001",  -- sqrt(1681) = 41
"000101001",  -- sqrt(1682) = 41
"000101001",  -- sqrt(1683) = 41
"000101001",  -- sqrt(1684) = 41
"000101001",  -- sqrt(1685) = 41
"000101001",  -- sqrt(1686) = 41
"000101001",  -- sqrt(1687) = 41
"000101001",  -- sqrt(1688) = 41
"000101001",  -- sqrt(1689) = 41
"000101001",  -- sqrt(1690) = 41
"000101001",  -- sqrt(1691) = 41
"000101001",  -- sqrt(1692) = 41
"000101001",  -- sqrt(1693) = 41
"000101001",  -- sqrt(1694) = 41
"000101001",  -- sqrt(1695) = 41
"000101001",  -- sqrt(1696) = 41
"000101001",  -- sqrt(1697) = 41
"000101001",  -- sqrt(1698) = 41
"000101001",  -- sqrt(1699) = 41
"000101001",  -- sqrt(1700) = 41
"000101001",  -- sqrt(1701) = 41
"000101001",  -- sqrt(1702) = 41
"000101001",  -- sqrt(1703) = 41
"000101001",  -- sqrt(1704) = 41
"000101001",  -- sqrt(1705) = 41
"000101001",  -- sqrt(1706) = 41
"000101001",  -- sqrt(1707) = 41
"000101001",  -- sqrt(1708) = 41
"000101001",  -- sqrt(1709) = 41
"000101001",  -- sqrt(1710) = 41
"000101001",  -- sqrt(1711) = 41
"000101001",  -- sqrt(1712) = 41
"000101001",  -- sqrt(1713) = 41
"000101001",  -- sqrt(1714) = 41
"000101001",  -- sqrt(1715) = 41
"000101001",  -- sqrt(1716) = 41
"000101001",  -- sqrt(1717) = 41
"000101001",  -- sqrt(1718) = 41
"000101001",  -- sqrt(1719) = 41
"000101001",  -- sqrt(1720) = 41
"000101001",  -- sqrt(1721) = 41
"000101001",  -- sqrt(1722) = 41
"000101010",  -- sqrt(1723) = 42
"000101010",  -- sqrt(1724) = 42
"000101010",  -- sqrt(1725) = 42
"000101010",  -- sqrt(1726) = 42
"000101010",  -- sqrt(1727) = 42
"000101010",  -- sqrt(1728) = 42
"000101010",  -- sqrt(1729) = 42
"000101010",  -- sqrt(1730) = 42
"000101010",  -- sqrt(1731) = 42
"000101010",  -- sqrt(1732) = 42
"000101010",  -- sqrt(1733) = 42
"000101010",  -- sqrt(1734) = 42
"000101010",  -- sqrt(1735) = 42
"000101010",  -- sqrt(1736) = 42
"000101010",  -- sqrt(1737) = 42
"000101010",  -- sqrt(1738) = 42
"000101010",  -- sqrt(1739) = 42
"000101010",  -- sqrt(1740) = 42
"000101010",  -- sqrt(1741) = 42
"000101010",  -- sqrt(1742) = 42
"000101010",  -- sqrt(1743) = 42
"000101010",  -- sqrt(1744) = 42
"000101010",  -- sqrt(1745) = 42
"000101010",  -- sqrt(1746) = 42
"000101010",  -- sqrt(1747) = 42
"000101010",  -- sqrt(1748) = 42
"000101010",  -- sqrt(1749) = 42
"000101010",  -- sqrt(1750) = 42
"000101010",  -- sqrt(1751) = 42
"000101010",  -- sqrt(1752) = 42
"000101010",  -- sqrt(1753) = 42
"000101010",  -- sqrt(1754) = 42
"000101010",  -- sqrt(1755) = 42
"000101010",  -- sqrt(1756) = 42
"000101010",  -- sqrt(1757) = 42
"000101010",  -- sqrt(1758) = 42
"000101010",  -- sqrt(1759) = 42
"000101010",  -- sqrt(1760) = 42
"000101010",  -- sqrt(1761) = 42
"000101010",  -- sqrt(1762) = 42
"000101010",  -- sqrt(1763) = 42
"000101010",  -- sqrt(1764) = 42
"000101010",  -- sqrt(1765) = 42
"000101010",  -- sqrt(1766) = 42
"000101010",  -- sqrt(1767) = 42
"000101010",  -- sqrt(1768) = 42
"000101010",  -- sqrt(1769) = 42
"000101010",  -- sqrt(1770) = 42
"000101010",  -- sqrt(1771) = 42
"000101010",  -- sqrt(1772) = 42
"000101010",  -- sqrt(1773) = 42
"000101010",  -- sqrt(1774) = 42
"000101010",  -- sqrt(1775) = 42
"000101010",  -- sqrt(1776) = 42
"000101010",  -- sqrt(1777) = 42
"000101010",  -- sqrt(1778) = 42
"000101010",  -- sqrt(1779) = 42
"000101010",  -- sqrt(1780) = 42
"000101010",  -- sqrt(1781) = 42
"000101010",  -- sqrt(1782) = 42
"000101010",  -- sqrt(1783) = 42
"000101010",  -- sqrt(1784) = 42
"000101010",  -- sqrt(1785) = 42
"000101010",  -- sqrt(1786) = 42
"000101010",  -- sqrt(1787) = 42
"000101010",  -- sqrt(1788) = 42
"000101010",  -- sqrt(1789) = 42
"000101010",  -- sqrt(1790) = 42
"000101010",  -- sqrt(1791) = 42
"000101010",  -- sqrt(1792) = 42
"000101010",  -- sqrt(1793) = 42
"000101010",  -- sqrt(1794) = 42
"000101010",  -- sqrt(1795) = 42
"000101010",  -- sqrt(1796) = 42
"000101010",  -- sqrt(1797) = 42
"000101010",  -- sqrt(1798) = 42
"000101010",  -- sqrt(1799) = 42
"000101010",  -- sqrt(1800) = 42
"000101010",  -- sqrt(1801) = 42
"000101010",  -- sqrt(1802) = 42
"000101010",  -- sqrt(1803) = 42
"000101010",  -- sqrt(1804) = 42
"000101010",  -- sqrt(1805) = 42
"000101010",  -- sqrt(1806) = 42
"000101011",  -- sqrt(1807) = 43
"000101011",  -- sqrt(1808) = 43
"000101011",  -- sqrt(1809) = 43
"000101011",  -- sqrt(1810) = 43
"000101011",  -- sqrt(1811) = 43
"000101011",  -- sqrt(1812) = 43
"000101011",  -- sqrt(1813) = 43
"000101011",  -- sqrt(1814) = 43
"000101011",  -- sqrt(1815) = 43
"000101011",  -- sqrt(1816) = 43
"000101011",  -- sqrt(1817) = 43
"000101011",  -- sqrt(1818) = 43
"000101011",  -- sqrt(1819) = 43
"000101011",  -- sqrt(1820) = 43
"000101011",  -- sqrt(1821) = 43
"000101011",  -- sqrt(1822) = 43
"000101011",  -- sqrt(1823) = 43
"000101011",  -- sqrt(1824) = 43
"000101011",  -- sqrt(1825) = 43
"000101011",  -- sqrt(1826) = 43
"000101011",  -- sqrt(1827) = 43
"000101011",  -- sqrt(1828) = 43
"000101011",  -- sqrt(1829) = 43
"000101011",  -- sqrt(1830) = 43
"000101011",  -- sqrt(1831) = 43
"000101011",  -- sqrt(1832) = 43
"000101011",  -- sqrt(1833) = 43
"000101011",  -- sqrt(1834) = 43
"000101011",  -- sqrt(1835) = 43
"000101011",  -- sqrt(1836) = 43
"000101011",  -- sqrt(1837) = 43
"000101011",  -- sqrt(1838) = 43
"000101011",  -- sqrt(1839) = 43
"000101011",  -- sqrt(1840) = 43
"000101011",  -- sqrt(1841) = 43
"000101011",  -- sqrt(1842) = 43
"000101011",  -- sqrt(1843) = 43
"000101011",  -- sqrt(1844) = 43
"000101011",  -- sqrt(1845) = 43
"000101011",  -- sqrt(1846) = 43
"000101011",  -- sqrt(1847) = 43
"000101011",  -- sqrt(1848) = 43
"000101011",  -- sqrt(1849) = 43
"000101011",  -- sqrt(1850) = 43
"000101011",  -- sqrt(1851) = 43
"000101011",  -- sqrt(1852) = 43
"000101011",  -- sqrt(1853) = 43
"000101011",  -- sqrt(1854) = 43
"000101011",  -- sqrt(1855) = 43
"000101011",  -- sqrt(1856) = 43
"000101011",  -- sqrt(1857) = 43
"000101011",  -- sqrt(1858) = 43
"000101011",  -- sqrt(1859) = 43
"000101011",  -- sqrt(1860) = 43
"000101011",  -- sqrt(1861) = 43
"000101011",  -- sqrt(1862) = 43
"000101011",  -- sqrt(1863) = 43
"000101011",  -- sqrt(1864) = 43
"000101011",  -- sqrt(1865) = 43
"000101011",  -- sqrt(1866) = 43
"000101011",  -- sqrt(1867) = 43
"000101011",  -- sqrt(1868) = 43
"000101011",  -- sqrt(1869) = 43
"000101011",  -- sqrt(1870) = 43
"000101011",  -- sqrt(1871) = 43
"000101011",  -- sqrt(1872) = 43
"000101011",  -- sqrt(1873) = 43
"000101011",  -- sqrt(1874) = 43
"000101011",  -- sqrt(1875) = 43
"000101011",  -- sqrt(1876) = 43
"000101011",  -- sqrt(1877) = 43
"000101011",  -- sqrt(1878) = 43
"000101011",  -- sqrt(1879) = 43
"000101011",  -- sqrt(1880) = 43
"000101011",  -- sqrt(1881) = 43
"000101011",  -- sqrt(1882) = 43
"000101011",  -- sqrt(1883) = 43
"000101011",  -- sqrt(1884) = 43
"000101011",  -- sqrt(1885) = 43
"000101011",  -- sqrt(1886) = 43
"000101011",  -- sqrt(1887) = 43
"000101011",  -- sqrt(1888) = 43
"000101011",  -- sqrt(1889) = 43
"000101011",  -- sqrt(1890) = 43
"000101011",  -- sqrt(1891) = 43
"000101011",  -- sqrt(1892) = 43
"000101100",  -- sqrt(1893) = 44
"000101100",  -- sqrt(1894) = 44
"000101100",  -- sqrt(1895) = 44
"000101100",  -- sqrt(1896) = 44
"000101100",  -- sqrt(1897) = 44
"000101100",  -- sqrt(1898) = 44
"000101100",  -- sqrt(1899) = 44
"000101100",  -- sqrt(1900) = 44
"000101100",  -- sqrt(1901) = 44
"000101100",  -- sqrt(1902) = 44
"000101100",  -- sqrt(1903) = 44
"000101100",  -- sqrt(1904) = 44
"000101100",  -- sqrt(1905) = 44
"000101100",  -- sqrt(1906) = 44
"000101100",  -- sqrt(1907) = 44
"000101100",  -- sqrt(1908) = 44
"000101100",  -- sqrt(1909) = 44
"000101100",  -- sqrt(1910) = 44
"000101100",  -- sqrt(1911) = 44
"000101100",  -- sqrt(1912) = 44
"000101100",  -- sqrt(1913) = 44
"000101100",  -- sqrt(1914) = 44
"000101100",  -- sqrt(1915) = 44
"000101100",  -- sqrt(1916) = 44
"000101100",  -- sqrt(1917) = 44
"000101100",  -- sqrt(1918) = 44
"000101100",  -- sqrt(1919) = 44
"000101100",  -- sqrt(1920) = 44
"000101100",  -- sqrt(1921) = 44
"000101100",  -- sqrt(1922) = 44
"000101100",  -- sqrt(1923) = 44
"000101100",  -- sqrt(1924) = 44
"000101100",  -- sqrt(1925) = 44
"000101100",  -- sqrt(1926) = 44
"000101100",  -- sqrt(1927) = 44
"000101100",  -- sqrt(1928) = 44
"000101100",  -- sqrt(1929) = 44
"000101100",  -- sqrt(1930) = 44
"000101100",  -- sqrt(1931) = 44
"000101100",  -- sqrt(1932) = 44
"000101100",  -- sqrt(1933) = 44
"000101100",  -- sqrt(1934) = 44
"000101100",  -- sqrt(1935) = 44
"000101100",  -- sqrt(1936) = 44
"000101100",  -- sqrt(1937) = 44
"000101100",  -- sqrt(1938) = 44
"000101100",  -- sqrt(1939) = 44
"000101100",  -- sqrt(1940) = 44
"000101100",  -- sqrt(1941) = 44
"000101100",  -- sqrt(1942) = 44
"000101100",  -- sqrt(1943) = 44
"000101100",  -- sqrt(1944) = 44
"000101100",  -- sqrt(1945) = 44
"000101100",  -- sqrt(1946) = 44
"000101100",  -- sqrt(1947) = 44
"000101100",  -- sqrt(1948) = 44
"000101100",  -- sqrt(1949) = 44
"000101100",  -- sqrt(1950) = 44
"000101100",  -- sqrt(1951) = 44
"000101100",  -- sqrt(1952) = 44
"000101100",  -- sqrt(1953) = 44
"000101100",  -- sqrt(1954) = 44
"000101100",  -- sqrt(1955) = 44
"000101100",  -- sqrt(1956) = 44
"000101100",  -- sqrt(1957) = 44
"000101100",  -- sqrt(1958) = 44
"000101100",  -- sqrt(1959) = 44
"000101100",  -- sqrt(1960) = 44
"000101100",  -- sqrt(1961) = 44
"000101100",  -- sqrt(1962) = 44
"000101100",  -- sqrt(1963) = 44
"000101100",  -- sqrt(1964) = 44
"000101100",  -- sqrt(1965) = 44
"000101100",  -- sqrt(1966) = 44
"000101100",  -- sqrt(1967) = 44
"000101100",  -- sqrt(1968) = 44
"000101100",  -- sqrt(1969) = 44
"000101100",  -- sqrt(1970) = 44
"000101100",  -- sqrt(1971) = 44
"000101100",  -- sqrt(1972) = 44
"000101100",  -- sqrt(1973) = 44
"000101100",  -- sqrt(1974) = 44
"000101100",  -- sqrt(1975) = 44
"000101100",  -- sqrt(1976) = 44
"000101100",  -- sqrt(1977) = 44
"000101100",  -- sqrt(1978) = 44
"000101100",  -- sqrt(1979) = 44
"000101100",  -- sqrt(1980) = 44
"000101101",  -- sqrt(1981) = 45
"000101101",  -- sqrt(1982) = 45
"000101101",  -- sqrt(1983) = 45
"000101101",  -- sqrt(1984) = 45
"000101101",  -- sqrt(1985) = 45
"000101101",  -- sqrt(1986) = 45
"000101101",  -- sqrt(1987) = 45
"000101101",  -- sqrt(1988) = 45
"000101101",  -- sqrt(1989) = 45
"000101101",  -- sqrt(1990) = 45
"000101101",  -- sqrt(1991) = 45
"000101101",  -- sqrt(1992) = 45
"000101101",  -- sqrt(1993) = 45
"000101101",  -- sqrt(1994) = 45
"000101101",  -- sqrt(1995) = 45
"000101101",  -- sqrt(1996) = 45
"000101101",  -- sqrt(1997) = 45
"000101101",  -- sqrt(1998) = 45
"000101101",  -- sqrt(1999) = 45
"000101101",  -- sqrt(2000) = 45
"000101101",  -- sqrt(2001) = 45
"000101101",  -- sqrt(2002) = 45
"000101101",  -- sqrt(2003) = 45
"000101101",  -- sqrt(2004) = 45
"000101101",  -- sqrt(2005) = 45
"000101101",  -- sqrt(2006) = 45
"000101101",  -- sqrt(2007) = 45
"000101101",  -- sqrt(2008) = 45
"000101101",  -- sqrt(2009) = 45
"000101101",  -- sqrt(2010) = 45
"000101101",  -- sqrt(2011) = 45
"000101101",  -- sqrt(2012) = 45
"000101101",  -- sqrt(2013) = 45
"000101101",  -- sqrt(2014) = 45
"000101101",  -- sqrt(2015) = 45
"000101101",  -- sqrt(2016) = 45
"000101101",  -- sqrt(2017) = 45
"000101101",  -- sqrt(2018) = 45
"000101101",  -- sqrt(2019) = 45
"000101101",  -- sqrt(2020) = 45
"000101101",  -- sqrt(2021) = 45
"000101101",  -- sqrt(2022) = 45
"000101101",  -- sqrt(2023) = 45
"000101101",  -- sqrt(2024) = 45
"000101101",  -- sqrt(2025) = 45
"000101101",  -- sqrt(2026) = 45
"000101101",  -- sqrt(2027) = 45
"000101101",  -- sqrt(2028) = 45
"000101101",  -- sqrt(2029) = 45
"000101101",  -- sqrt(2030) = 45
"000101101",  -- sqrt(2031) = 45
"000101101",  -- sqrt(2032) = 45
"000101101",  -- sqrt(2033) = 45
"000101101",  -- sqrt(2034) = 45
"000101101",  -- sqrt(2035) = 45
"000101101",  -- sqrt(2036) = 45
"000101101",  -- sqrt(2037) = 45
"000101101",  -- sqrt(2038) = 45
"000101101",  -- sqrt(2039) = 45
"000101101",  -- sqrt(2040) = 45
"000101101",  -- sqrt(2041) = 45
"000101101",  -- sqrt(2042) = 45
"000101101",  -- sqrt(2043) = 45
"000101101",  -- sqrt(2044) = 45
"000101101",  -- sqrt(2045) = 45
"000101101",  -- sqrt(2046) = 45
"000101101",  -- sqrt(2047) = 45
"000101101",  -- sqrt(2048) = 45
"000101101",  -- sqrt(2049) = 45
"000101101",  -- sqrt(2050) = 45
"000101101",  -- sqrt(2051) = 45
"000101101",  -- sqrt(2052) = 45
"000101101",  -- sqrt(2053) = 45
"000101101",  -- sqrt(2054) = 45
"000101101",  -- sqrt(2055) = 45
"000101101",  -- sqrt(2056) = 45
"000101101",  -- sqrt(2057) = 45
"000101101",  -- sqrt(2058) = 45
"000101101",  -- sqrt(2059) = 45
"000101101",  -- sqrt(2060) = 45
"000101101",  -- sqrt(2061) = 45
"000101101",  -- sqrt(2062) = 45
"000101101",  -- sqrt(2063) = 45
"000101101",  -- sqrt(2064) = 45
"000101101",  -- sqrt(2065) = 45
"000101101",  -- sqrt(2066) = 45
"000101101",  -- sqrt(2067) = 45
"000101101",  -- sqrt(2068) = 45
"000101101",  -- sqrt(2069) = 45
"000101101",  -- sqrt(2070) = 45
"000101110",  -- sqrt(2071) = 46
"000101110",  -- sqrt(2072) = 46
"000101110",  -- sqrt(2073) = 46
"000101110",  -- sqrt(2074) = 46
"000101110",  -- sqrt(2075) = 46
"000101110",  -- sqrt(2076) = 46
"000101110",  -- sqrt(2077) = 46
"000101110",  -- sqrt(2078) = 46
"000101110",  -- sqrt(2079) = 46
"000101110",  -- sqrt(2080) = 46
"000101110",  -- sqrt(2081) = 46
"000101110",  -- sqrt(2082) = 46
"000101110",  -- sqrt(2083) = 46
"000101110",  -- sqrt(2084) = 46
"000101110",  -- sqrt(2085) = 46
"000101110",  -- sqrt(2086) = 46
"000101110",  -- sqrt(2087) = 46
"000101110",  -- sqrt(2088) = 46
"000101110",  -- sqrt(2089) = 46
"000101110",  -- sqrt(2090) = 46
"000101110",  -- sqrt(2091) = 46
"000101110",  -- sqrt(2092) = 46
"000101110",  -- sqrt(2093) = 46
"000101110",  -- sqrt(2094) = 46
"000101110",  -- sqrt(2095) = 46
"000101110",  -- sqrt(2096) = 46
"000101110",  -- sqrt(2097) = 46
"000101110",  -- sqrt(2098) = 46
"000101110",  -- sqrt(2099) = 46
"000101110",  -- sqrt(2100) = 46
"000101110",  -- sqrt(2101) = 46
"000101110",  -- sqrt(2102) = 46
"000101110",  -- sqrt(2103) = 46
"000101110",  -- sqrt(2104) = 46
"000101110",  -- sqrt(2105) = 46
"000101110",  -- sqrt(2106) = 46
"000101110",  -- sqrt(2107) = 46
"000101110",  -- sqrt(2108) = 46
"000101110",  -- sqrt(2109) = 46
"000101110",  -- sqrt(2110) = 46
"000101110",  -- sqrt(2111) = 46
"000101110",  -- sqrt(2112) = 46
"000101110",  -- sqrt(2113) = 46
"000101110",  -- sqrt(2114) = 46
"000101110",  -- sqrt(2115) = 46
"000101110",  -- sqrt(2116) = 46
"000101110",  -- sqrt(2117) = 46
"000101110",  -- sqrt(2118) = 46
"000101110",  -- sqrt(2119) = 46
"000101110",  -- sqrt(2120) = 46
"000101110",  -- sqrt(2121) = 46
"000101110",  -- sqrt(2122) = 46
"000101110",  -- sqrt(2123) = 46
"000101110",  -- sqrt(2124) = 46
"000101110",  -- sqrt(2125) = 46
"000101110",  -- sqrt(2126) = 46
"000101110",  -- sqrt(2127) = 46
"000101110",  -- sqrt(2128) = 46
"000101110",  -- sqrt(2129) = 46
"000101110",  -- sqrt(2130) = 46
"000101110",  -- sqrt(2131) = 46
"000101110",  -- sqrt(2132) = 46
"000101110",  -- sqrt(2133) = 46
"000101110",  -- sqrt(2134) = 46
"000101110",  -- sqrt(2135) = 46
"000101110",  -- sqrt(2136) = 46
"000101110",  -- sqrt(2137) = 46
"000101110",  -- sqrt(2138) = 46
"000101110",  -- sqrt(2139) = 46
"000101110",  -- sqrt(2140) = 46
"000101110",  -- sqrt(2141) = 46
"000101110",  -- sqrt(2142) = 46
"000101110",  -- sqrt(2143) = 46
"000101110",  -- sqrt(2144) = 46
"000101110",  -- sqrt(2145) = 46
"000101110",  -- sqrt(2146) = 46
"000101110",  -- sqrt(2147) = 46
"000101110",  -- sqrt(2148) = 46
"000101110",  -- sqrt(2149) = 46
"000101110",  -- sqrt(2150) = 46
"000101110",  -- sqrt(2151) = 46
"000101110",  -- sqrt(2152) = 46
"000101110",  -- sqrt(2153) = 46
"000101110",  -- sqrt(2154) = 46
"000101110",  -- sqrt(2155) = 46
"000101110",  -- sqrt(2156) = 46
"000101110",  -- sqrt(2157) = 46
"000101110",  -- sqrt(2158) = 46
"000101110",  -- sqrt(2159) = 46
"000101110",  -- sqrt(2160) = 46
"000101110",  -- sqrt(2161) = 46
"000101110",  -- sqrt(2162) = 46
"000101111",  -- sqrt(2163) = 47
"000101111",  -- sqrt(2164) = 47
"000101111",  -- sqrt(2165) = 47
"000101111",  -- sqrt(2166) = 47
"000101111",  -- sqrt(2167) = 47
"000101111",  -- sqrt(2168) = 47
"000101111",  -- sqrt(2169) = 47
"000101111",  -- sqrt(2170) = 47
"000101111",  -- sqrt(2171) = 47
"000101111",  -- sqrt(2172) = 47
"000101111",  -- sqrt(2173) = 47
"000101111",  -- sqrt(2174) = 47
"000101111",  -- sqrt(2175) = 47
"000101111",  -- sqrt(2176) = 47
"000101111",  -- sqrt(2177) = 47
"000101111",  -- sqrt(2178) = 47
"000101111",  -- sqrt(2179) = 47
"000101111",  -- sqrt(2180) = 47
"000101111",  -- sqrt(2181) = 47
"000101111",  -- sqrt(2182) = 47
"000101111",  -- sqrt(2183) = 47
"000101111",  -- sqrt(2184) = 47
"000101111",  -- sqrt(2185) = 47
"000101111",  -- sqrt(2186) = 47
"000101111",  -- sqrt(2187) = 47
"000101111",  -- sqrt(2188) = 47
"000101111",  -- sqrt(2189) = 47
"000101111",  -- sqrt(2190) = 47
"000101111",  -- sqrt(2191) = 47
"000101111",  -- sqrt(2192) = 47
"000101111",  -- sqrt(2193) = 47
"000101111",  -- sqrt(2194) = 47
"000101111",  -- sqrt(2195) = 47
"000101111",  -- sqrt(2196) = 47
"000101111",  -- sqrt(2197) = 47
"000101111",  -- sqrt(2198) = 47
"000101111",  -- sqrt(2199) = 47
"000101111",  -- sqrt(2200) = 47
"000101111",  -- sqrt(2201) = 47
"000101111",  -- sqrt(2202) = 47
"000101111",  -- sqrt(2203) = 47
"000101111",  -- sqrt(2204) = 47
"000101111",  -- sqrt(2205) = 47
"000101111",  -- sqrt(2206) = 47
"000101111",  -- sqrt(2207) = 47
"000101111",  -- sqrt(2208) = 47
"000101111",  -- sqrt(2209) = 47
"000101111",  -- sqrt(2210) = 47
"000101111",  -- sqrt(2211) = 47
"000101111",  -- sqrt(2212) = 47
"000101111",  -- sqrt(2213) = 47
"000101111",  -- sqrt(2214) = 47
"000101111",  -- sqrt(2215) = 47
"000101111",  -- sqrt(2216) = 47
"000101111",  -- sqrt(2217) = 47
"000101111",  -- sqrt(2218) = 47
"000101111",  -- sqrt(2219) = 47
"000101111",  -- sqrt(2220) = 47
"000101111",  -- sqrt(2221) = 47
"000101111",  -- sqrt(2222) = 47
"000101111",  -- sqrt(2223) = 47
"000101111",  -- sqrt(2224) = 47
"000101111",  -- sqrt(2225) = 47
"000101111",  -- sqrt(2226) = 47
"000101111",  -- sqrt(2227) = 47
"000101111",  -- sqrt(2228) = 47
"000101111",  -- sqrt(2229) = 47
"000101111",  -- sqrt(2230) = 47
"000101111",  -- sqrt(2231) = 47
"000101111",  -- sqrt(2232) = 47
"000101111",  -- sqrt(2233) = 47
"000101111",  -- sqrt(2234) = 47
"000101111",  -- sqrt(2235) = 47
"000101111",  -- sqrt(2236) = 47
"000101111",  -- sqrt(2237) = 47
"000101111",  -- sqrt(2238) = 47
"000101111",  -- sqrt(2239) = 47
"000101111",  -- sqrt(2240) = 47
"000101111",  -- sqrt(2241) = 47
"000101111",  -- sqrt(2242) = 47
"000101111",  -- sqrt(2243) = 47
"000101111",  -- sqrt(2244) = 47
"000101111",  -- sqrt(2245) = 47
"000101111",  -- sqrt(2246) = 47
"000101111",  -- sqrt(2247) = 47
"000101111",  -- sqrt(2248) = 47
"000101111",  -- sqrt(2249) = 47
"000101111",  -- sqrt(2250) = 47
"000101111",  -- sqrt(2251) = 47
"000101111",  -- sqrt(2252) = 47
"000101111",  -- sqrt(2253) = 47
"000101111",  -- sqrt(2254) = 47
"000101111",  -- sqrt(2255) = 47
"000101111",  -- sqrt(2256) = 47
"000110000",  -- sqrt(2257) = 48
"000110000",  -- sqrt(2258) = 48
"000110000",  -- sqrt(2259) = 48
"000110000",  -- sqrt(2260) = 48
"000110000",  -- sqrt(2261) = 48
"000110000",  -- sqrt(2262) = 48
"000110000",  -- sqrt(2263) = 48
"000110000",  -- sqrt(2264) = 48
"000110000",  -- sqrt(2265) = 48
"000110000",  -- sqrt(2266) = 48
"000110000",  -- sqrt(2267) = 48
"000110000",  -- sqrt(2268) = 48
"000110000",  -- sqrt(2269) = 48
"000110000",  -- sqrt(2270) = 48
"000110000",  -- sqrt(2271) = 48
"000110000",  -- sqrt(2272) = 48
"000110000",  -- sqrt(2273) = 48
"000110000",  -- sqrt(2274) = 48
"000110000",  -- sqrt(2275) = 48
"000110000",  -- sqrt(2276) = 48
"000110000",  -- sqrt(2277) = 48
"000110000",  -- sqrt(2278) = 48
"000110000",  -- sqrt(2279) = 48
"000110000",  -- sqrt(2280) = 48
"000110000",  -- sqrt(2281) = 48
"000110000",  -- sqrt(2282) = 48
"000110000",  -- sqrt(2283) = 48
"000110000",  -- sqrt(2284) = 48
"000110000",  -- sqrt(2285) = 48
"000110000",  -- sqrt(2286) = 48
"000110000",  -- sqrt(2287) = 48
"000110000",  -- sqrt(2288) = 48
"000110000",  -- sqrt(2289) = 48
"000110000",  -- sqrt(2290) = 48
"000110000",  -- sqrt(2291) = 48
"000110000",  -- sqrt(2292) = 48
"000110000",  -- sqrt(2293) = 48
"000110000",  -- sqrt(2294) = 48
"000110000",  -- sqrt(2295) = 48
"000110000",  -- sqrt(2296) = 48
"000110000",  -- sqrt(2297) = 48
"000110000",  -- sqrt(2298) = 48
"000110000",  -- sqrt(2299) = 48
"000110000",  -- sqrt(2300) = 48
"000110000",  -- sqrt(2301) = 48
"000110000",  -- sqrt(2302) = 48
"000110000",  -- sqrt(2303) = 48
"000110000",  -- sqrt(2304) = 48
"000110000",  -- sqrt(2305) = 48
"000110000",  -- sqrt(2306) = 48
"000110000",  -- sqrt(2307) = 48
"000110000",  -- sqrt(2308) = 48
"000110000",  -- sqrt(2309) = 48
"000110000",  -- sqrt(2310) = 48
"000110000",  -- sqrt(2311) = 48
"000110000",  -- sqrt(2312) = 48
"000110000",  -- sqrt(2313) = 48
"000110000",  -- sqrt(2314) = 48
"000110000",  -- sqrt(2315) = 48
"000110000",  -- sqrt(2316) = 48
"000110000",  -- sqrt(2317) = 48
"000110000",  -- sqrt(2318) = 48
"000110000",  -- sqrt(2319) = 48
"000110000",  -- sqrt(2320) = 48
"000110000",  -- sqrt(2321) = 48
"000110000",  -- sqrt(2322) = 48
"000110000",  -- sqrt(2323) = 48
"000110000",  -- sqrt(2324) = 48
"000110000",  -- sqrt(2325) = 48
"000110000",  -- sqrt(2326) = 48
"000110000",  -- sqrt(2327) = 48
"000110000",  -- sqrt(2328) = 48
"000110000",  -- sqrt(2329) = 48
"000110000",  -- sqrt(2330) = 48
"000110000",  -- sqrt(2331) = 48
"000110000",  -- sqrt(2332) = 48
"000110000",  -- sqrt(2333) = 48
"000110000",  -- sqrt(2334) = 48
"000110000",  -- sqrt(2335) = 48
"000110000",  -- sqrt(2336) = 48
"000110000",  -- sqrt(2337) = 48
"000110000",  -- sqrt(2338) = 48
"000110000",  -- sqrt(2339) = 48
"000110000",  -- sqrt(2340) = 48
"000110000",  -- sqrt(2341) = 48
"000110000",  -- sqrt(2342) = 48
"000110000",  -- sqrt(2343) = 48
"000110000",  -- sqrt(2344) = 48
"000110000",  -- sqrt(2345) = 48
"000110000",  -- sqrt(2346) = 48
"000110000",  -- sqrt(2347) = 48
"000110000",  -- sqrt(2348) = 48
"000110000",  -- sqrt(2349) = 48
"000110000",  -- sqrt(2350) = 48
"000110000",  -- sqrt(2351) = 48
"000110000",  -- sqrt(2352) = 48
"000110001",  -- sqrt(2353) = 49
"000110001",  -- sqrt(2354) = 49
"000110001",  -- sqrt(2355) = 49
"000110001",  -- sqrt(2356) = 49
"000110001",  -- sqrt(2357) = 49
"000110001",  -- sqrt(2358) = 49
"000110001",  -- sqrt(2359) = 49
"000110001",  -- sqrt(2360) = 49
"000110001",  -- sqrt(2361) = 49
"000110001",  -- sqrt(2362) = 49
"000110001",  -- sqrt(2363) = 49
"000110001",  -- sqrt(2364) = 49
"000110001",  -- sqrt(2365) = 49
"000110001",  -- sqrt(2366) = 49
"000110001",  -- sqrt(2367) = 49
"000110001",  -- sqrt(2368) = 49
"000110001",  -- sqrt(2369) = 49
"000110001",  -- sqrt(2370) = 49
"000110001",  -- sqrt(2371) = 49
"000110001",  -- sqrt(2372) = 49
"000110001",  -- sqrt(2373) = 49
"000110001",  -- sqrt(2374) = 49
"000110001",  -- sqrt(2375) = 49
"000110001",  -- sqrt(2376) = 49
"000110001",  -- sqrt(2377) = 49
"000110001",  -- sqrt(2378) = 49
"000110001",  -- sqrt(2379) = 49
"000110001",  -- sqrt(2380) = 49
"000110001",  -- sqrt(2381) = 49
"000110001",  -- sqrt(2382) = 49
"000110001",  -- sqrt(2383) = 49
"000110001",  -- sqrt(2384) = 49
"000110001",  -- sqrt(2385) = 49
"000110001",  -- sqrt(2386) = 49
"000110001",  -- sqrt(2387) = 49
"000110001",  -- sqrt(2388) = 49
"000110001",  -- sqrt(2389) = 49
"000110001",  -- sqrt(2390) = 49
"000110001",  -- sqrt(2391) = 49
"000110001",  -- sqrt(2392) = 49
"000110001",  -- sqrt(2393) = 49
"000110001",  -- sqrt(2394) = 49
"000110001",  -- sqrt(2395) = 49
"000110001",  -- sqrt(2396) = 49
"000110001",  -- sqrt(2397) = 49
"000110001",  -- sqrt(2398) = 49
"000110001",  -- sqrt(2399) = 49
"000110001",  -- sqrt(2400) = 49
"000110001",  -- sqrt(2401) = 49
"000110001",  -- sqrt(2402) = 49
"000110001",  -- sqrt(2403) = 49
"000110001",  -- sqrt(2404) = 49
"000110001",  -- sqrt(2405) = 49
"000110001",  -- sqrt(2406) = 49
"000110001",  -- sqrt(2407) = 49
"000110001",  -- sqrt(2408) = 49
"000110001",  -- sqrt(2409) = 49
"000110001",  -- sqrt(2410) = 49
"000110001",  -- sqrt(2411) = 49
"000110001",  -- sqrt(2412) = 49
"000110001",  -- sqrt(2413) = 49
"000110001",  -- sqrt(2414) = 49
"000110001",  -- sqrt(2415) = 49
"000110001",  -- sqrt(2416) = 49
"000110001",  -- sqrt(2417) = 49
"000110001",  -- sqrt(2418) = 49
"000110001",  -- sqrt(2419) = 49
"000110001",  -- sqrt(2420) = 49
"000110001",  -- sqrt(2421) = 49
"000110001",  -- sqrt(2422) = 49
"000110001",  -- sqrt(2423) = 49
"000110001",  -- sqrt(2424) = 49
"000110001",  -- sqrt(2425) = 49
"000110001",  -- sqrt(2426) = 49
"000110001",  -- sqrt(2427) = 49
"000110001",  -- sqrt(2428) = 49
"000110001",  -- sqrt(2429) = 49
"000110001",  -- sqrt(2430) = 49
"000110001",  -- sqrt(2431) = 49
"000110001",  -- sqrt(2432) = 49
"000110001",  -- sqrt(2433) = 49
"000110001",  -- sqrt(2434) = 49
"000110001",  -- sqrt(2435) = 49
"000110001",  -- sqrt(2436) = 49
"000110001",  -- sqrt(2437) = 49
"000110001",  -- sqrt(2438) = 49
"000110001",  -- sqrt(2439) = 49
"000110001",  -- sqrt(2440) = 49
"000110001",  -- sqrt(2441) = 49
"000110001",  -- sqrt(2442) = 49
"000110001",  -- sqrt(2443) = 49
"000110001",  -- sqrt(2444) = 49
"000110001",  -- sqrt(2445) = 49
"000110001",  -- sqrt(2446) = 49
"000110001",  -- sqrt(2447) = 49
"000110001",  -- sqrt(2448) = 49
"000110001",  -- sqrt(2449) = 49
"000110001",  -- sqrt(2450) = 49
"000110010",  -- sqrt(2451) = 50
"000110010",  -- sqrt(2452) = 50
"000110010",  -- sqrt(2453) = 50
"000110010",  -- sqrt(2454) = 50
"000110010",  -- sqrt(2455) = 50
"000110010",  -- sqrt(2456) = 50
"000110010",  -- sqrt(2457) = 50
"000110010",  -- sqrt(2458) = 50
"000110010",  -- sqrt(2459) = 50
"000110010",  -- sqrt(2460) = 50
"000110010",  -- sqrt(2461) = 50
"000110010",  -- sqrt(2462) = 50
"000110010",  -- sqrt(2463) = 50
"000110010",  -- sqrt(2464) = 50
"000110010",  -- sqrt(2465) = 50
"000110010",  -- sqrt(2466) = 50
"000110010",  -- sqrt(2467) = 50
"000110010",  -- sqrt(2468) = 50
"000110010",  -- sqrt(2469) = 50
"000110010",  -- sqrt(2470) = 50
"000110010",  -- sqrt(2471) = 50
"000110010",  -- sqrt(2472) = 50
"000110010",  -- sqrt(2473) = 50
"000110010",  -- sqrt(2474) = 50
"000110010",  -- sqrt(2475) = 50
"000110010",  -- sqrt(2476) = 50
"000110010",  -- sqrt(2477) = 50
"000110010",  -- sqrt(2478) = 50
"000110010",  -- sqrt(2479) = 50
"000110010",  -- sqrt(2480) = 50
"000110010",  -- sqrt(2481) = 50
"000110010",  -- sqrt(2482) = 50
"000110010",  -- sqrt(2483) = 50
"000110010",  -- sqrt(2484) = 50
"000110010",  -- sqrt(2485) = 50
"000110010",  -- sqrt(2486) = 50
"000110010",  -- sqrt(2487) = 50
"000110010",  -- sqrt(2488) = 50
"000110010",  -- sqrt(2489) = 50
"000110010",  -- sqrt(2490) = 50
"000110010",  -- sqrt(2491) = 50
"000110010",  -- sqrt(2492) = 50
"000110010",  -- sqrt(2493) = 50
"000110010",  -- sqrt(2494) = 50
"000110010",  -- sqrt(2495) = 50
"000110010",  -- sqrt(2496) = 50
"000110010",  -- sqrt(2497) = 50
"000110010",  -- sqrt(2498) = 50
"000110010",  -- sqrt(2499) = 50
"000110010",  -- sqrt(2500) = 50
"000110010",  -- sqrt(2501) = 50
"000110010",  -- sqrt(2502) = 50
"000110010",  -- sqrt(2503) = 50
"000110010",  -- sqrt(2504) = 50
"000110010",  -- sqrt(2505) = 50
"000110010",  -- sqrt(2506) = 50
"000110010",  -- sqrt(2507) = 50
"000110010",  -- sqrt(2508) = 50
"000110010",  -- sqrt(2509) = 50
"000110010",  -- sqrt(2510) = 50
"000110010",  -- sqrt(2511) = 50
"000110010",  -- sqrt(2512) = 50
"000110010",  -- sqrt(2513) = 50
"000110010",  -- sqrt(2514) = 50
"000110010",  -- sqrt(2515) = 50
"000110010",  -- sqrt(2516) = 50
"000110010",  -- sqrt(2517) = 50
"000110010",  -- sqrt(2518) = 50
"000110010",  -- sqrt(2519) = 50
"000110010",  -- sqrt(2520) = 50
"000110010",  -- sqrt(2521) = 50
"000110010",  -- sqrt(2522) = 50
"000110010",  -- sqrt(2523) = 50
"000110010",  -- sqrt(2524) = 50
"000110010",  -- sqrt(2525) = 50
"000110010",  -- sqrt(2526) = 50
"000110010",  -- sqrt(2527) = 50
"000110010",  -- sqrt(2528) = 50
"000110010",  -- sqrt(2529) = 50
"000110010",  -- sqrt(2530) = 50
"000110010",  -- sqrt(2531) = 50
"000110010",  -- sqrt(2532) = 50
"000110010",  -- sqrt(2533) = 50
"000110010",  -- sqrt(2534) = 50
"000110010",  -- sqrt(2535) = 50
"000110010",  -- sqrt(2536) = 50
"000110010",  -- sqrt(2537) = 50
"000110010",  -- sqrt(2538) = 50
"000110010",  -- sqrt(2539) = 50
"000110010",  -- sqrt(2540) = 50
"000110010",  -- sqrt(2541) = 50
"000110010",  -- sqrt(2542) = 50
"000110010",  -- sqrt(2543) = 50
"000110010",  -- sqrt(2544) = 50
"000110010",  -- sqrt(2545) = 50
"000110010",  -- sqrt(2546) = 50
"000110010",  -- sqrt(2547) = 50
"000110010",  -- sqrt(2548) = 50
"000110010",  -- sqrt(2549) = 50
"000110010",  -- sqrt(2550) = 50
"000110011",  -- sqrt(2551) = 51
"000110011",  -- sqrt(2552) = 51
"000110011",  -- sqrt(2553) = 51
"000110011",  -- sqrt(2554) = 51
"000110011",  -- sqrt(2555) = 51
"000110011",  -- sqrt(2556) = 51
"000110011",  -- sqrt(2557) = 51
"000110011",  -- sqrt(2558) = 51
"000110011",  -- sqrt(2559) = 51
"000110011",  -- sqrt(2560) = 51
"000110011",  -- sqrt(2561) = 51
"000110011",  -- sqrt(2562) = 51
"000110011",  -- sqrt(2563) = 51
"000110011",  -- sqrt(2564) = 51
"000110011",  -- sqrt(2565) = 51
"000110011",  -- sqrt(2566) = 51
"000110011",  -- sqrt(2567) = 51
"000110011",  -- sqrt(2568) = 51
"000110011",  -- sqrt(2569) = 51
"000110011",  -- sqrt(2570) = 51
"000110011",  -- sqrt(2571) = 51
"000110011",  -- sqrt(2572) = 51
"000110011",  -- sqrt(2573) = 51
"000110011",  -- sqrt(2574) = 51
"000110011",  -- sqrt(2575) = 51
"000110011",  -- sqrt(2576) = 51
"000110011",  -- sqrt(2577) = 51
"000110011",  -- sqrt(2578) = 51
"000110011",  -- sqrt(2579) = 51
"000110011",  -- sqrt(2580) = 51
"000110011",  -- sqrt(2581) = 51
"000110011",  -- sqrt(2582) = 51
"000110011",  -- sqrt(2583) = 51
"000110011",  -- sqrt(2584) = 51
"000110011",  -- sqrt(2585) = 51
"000110011",  -- sqrt(2586) = 51
"000110011",  -- sqrt(2587) = 51
"000110011",  -- sqrt(2588) = 51
"000110011",  -- sqrt(2589) = 51
"000110011",  -- sqrt(2590) = 51
"000110011",  -- sqrt(2591) = 51
"000110011",  -- sqrt(2592) = 51
"000110011",  -- sqrt(2593) = 51
"000110011",  -- sqrt(2594) = 51
"000110011",  -- sqrt(2595) = 51
"000110011",  -- sqrt(2596) = 51
"000110011",  -- sqrt(2597) = 51
"000110011",  -- sqrt(2598) = 51
"000110011",  -- sqrt(2599) = 51
"000110011",  -- sqrt(2600) = 51
"000110011",  -- sqrt(2601) = 51
"000110011",  -- sqrt(2602) = 51
"000110011",  -- sqrt(2603) = 51
"000110011",  -- sqrt(2604) = 51
"000110011",  -- sqrt(2605) = 51
"000110011",  -- sqrt(2606) = 51
"000110011",  -- sqrt(2607) = 51
"000110011",  -- sqrt(2608) = 51
"000110011",  -- sqrt(2609) = 51
"000110011",  -- sqrt(2610) = 51
"000110011",  -- sqrt(2611) = 51
"000110011",  -- sqrt(2612) = 51
"000110011",  -- sqrt(2613) = 51
"000110011",  -- sqrt(2614) = 51
"000110011",  -- sqrt(2615) = 51
"000110011",  -- sqrt(2616) = 51
"000110011",  -- sqrt(2617) = 51
"000110011",  -- sqrt(2618) = 51
"000110011",  -- sqrt(2619) = 51
"000110011",  -- sqrt(2620) = 51
"000110011",  -- sqrt(2621) = 51
"000110011",  -- sqrt(2622) = 51
"000110011",  -- sqrt(2623) = 51
"000110011",  -- sqrt(2624) = 51
"000110011",  -- sqrt(2625) = 51
"000110011",  -- sqrt(2626) = 51
"000110011",  -- sqrt(2627) = 51
"000110011",  -- sqrt(2628) = 51
"000110011",  -- sqrt(2629) = 51
"000110011",  -- sqrt(2630) = 51
"000110011",  -- sqrt(2631) = 51
"000110011",  -- sqrt(2632) = 51
"000110011",  -- sqrt(2633) = 51
"000110011",  -- sqrt(2634) = 51
"000110011",  -- sqrt(2635) = 51
"000110011",  -- sqrt(2636) = 51
"000110011",  -- sqrt(2637) = 51
"000110011",  -- sqrt(2638) = 51
"000110011",  -- sqrt(2639) = 51
"000110011",  -- sqrt(2640) = 51
"000110011",  -- sqrt(2641) = 51
"000110011",  -- sqrt(2642) = 51
"000110011",  -- sqrt(2643) = 51
"000110011",  -- sqrt(2644) = 51
"000110011",  -- sqrt(2645) = 51
"000110011",  -- sqrt(2646) = 51
"000110011",  -- sqrt(2647) = 51
"000110011",  -- sqrt(2648) = 51
"000110011",  -- sqrt(2649) = 51
"000110011",  -- sqrt(2650) = 51
"000110011",  -- sqrt(2651) = 51
"000110011",  -- sqrt(2652) = 51
"000110100",  -- sqrt(2653) = 52
"000110100",  -- sqrt(2654) = 52
"000110100",  -- sqrt(2655) = 52
"000110100",  -- sqrt(2656) = 52
"000110100",  -- sqrt(2657) = 52
"000110100",  -- sqrt(2658) = 52
"000110100",  -- sqrt(2659) = 52
"000110100",  -- sqrt(2660) = 52
"000110100",  -- sqrt(2661) = 52
"000110100",  -- sqrt(2662) = 52
"000110100",  -- sqrt(2663) = 52
"000110100",  -- sqrt(2664) = 52
"000110100",  -- sqrt(2665) = 52
"000110100",  -- sqrt(2666) = 52
"000110100",  -- sqrt(2667) = 52
"000110100",  -- sqrt(2668) = 52
"000110100",  -- sqrt(2669) = 52
"000110100",  -- sqrt(2670) = 52
"000110100",  -- sqrt(2671) = 52
"000110100",  -- sqrt(2672) = 52
"000110100",  -- sqrt(2673) = 52
"000110100",  -- sqrt(2674) = 52
"000110100",  -- sqrt(2675) = 52
"000110100",  -- sqrt(2676) = 52
"000110100",  -- sqrt(2677) = 52
"000110100",  -- sqrt(2678) = 52
"000110100",  -- sqrt(2679) = 52
"000110100",  -- sqrt(2680) = 52
"000110100",  -- sqrt(2681) = 52
"000110100",  -- sqrt(2682) = 52
"000110100",  -- sqrt(2683) = 52
"000110100",  -- sqrt(2684) = 52
"000110100",  -- sqrt(2685) = 52
"000110100",  -- sqrt(2686) = 52
"000110100",  -- sqrt(2687) = 52
"000110100",  -- sqrt(2688) = 52
"000110100",  -- sqrt(2689) = 52
"000110100",  -- sqrt(2690) = 52
"000110100",  -- sqrt(2691) = 52
"000110100",  -- sqrt(2692) = 52
"000110100",  -- sqrt(2693) = 52
"000110100",  -- sqrt(2694) = 52
"000110100",  -- sqrt(2695) = 52
"000110100",  -- sqrt(2696) = 52
"000110100",  -- sqrt(2697) = 52
"000110100",  -- sqrt(2698) = 52
"000110100",  -- sqrt(2699) = 52
"000110100",  -- sqrt(2700) = 52
"000110100",  -- sqrt(2701) = 52
"000110100",  -- sqrt(2702) = 52
"000110100",  -- sqrt(2703) = 52
"000110100",  -- sqrt(2704) = 52
"000110100",  -- sqrt(2705) = 52
"000110100",  -- sqrt(2706) = 52
"000110100",  -- sqrt(2707) = 52
"000110100",  -- sqrt(2708) = 52
"000110100",  -- sqrt(2709) = 52
"000110100",  -- sqrt(2710) = 52
"000110100",  -- sqrt(2711) = 52
"000110100",  -- sqrt(2712) = 52
"000110100",  -- sqrt(2713) = 52
"000110100",  -- sqrt(2714) = 52
"000110100",  -- sqrt(2715) = 52
"000110100",  -- sqrt(2716) = 52
"000110100",  -- sqrt(2717) = 52
"000110100",  -- sqrt(2718) = 52
"000110100",  -- sqrt(2719) = 52
"000110100",  -- sqrt(2720) = 52
"000110100",  -- sqrt(2721) = 52
"000110100",  -- sqrt(2722) = 52
"000110100",  -- sqrt(2723) = 52
"000110100",  -- sqrt(2724) = 52
"000110100",  -- sqrt(2725) = 52
"000110100",  -- sqrt(2726) = 52
"000110100",  -- sqrt(2727) = 52
"000110100",  -- sqrt(2728) = 52
"000110100",  -- sqrt(2729) = 52
"000110100",  -- sqrt(2730) = 52
"000110100",  -- sqrt(2731) = 52
"000110100",  -- sqrt(2732) = 52
"000110100",  -- sqrt(2733) = 52
"000110100",  -- sqrt(2734) = 52
"000110100",  -- sqrt(2735) = 52
"000110100",  -- sqrt(2736) = 52
"000110100",  -- sqrt(2737) = 52
"000110100",  -- sqrt(2738) = 52
"000110100",  -- sqrt(2739) = 52
"000110100",  -- sqrt(2740) = 52
"000110100",  -- sqrt(2741) = 52
"000110100",  -- sqrt(2742) = 52
"000110100",  -- sqrt(2743) = 52
"000110100",  -- sqrt(2744) = 52
"000110100",  -- sqrt(2745) = 52
"000110100",  -- sqrt(2746) = 52
"000110100",  -- sqrt(2747) = 52
"000110100",  -- sqrt(2748) = 52
"000110100",  -- sqrt(2749) = 52
"000110100",  -- sqrt(2750) = 52
"000110100",  -- sqrt(2751) = 52
"000110100",  -- sqrt(2752) = 52
"000110100",  -- sqrt(2753) = 52
"000110100",  -- sqrt(2754) = 52
"000110100",  -- sqrt(2755) = 52
"000110100",  -- sqrt(2756) = 52
"000110101",  -- sqrt(2757) = 53
"000110101",  -- sqrt(2758) = 53
"000110101",  -- sqrt(2759) = 53
"000110101",  -- sqrt(2760) = 53
"000110101",  -- sqrt(2761) = 53
"000110101",  -- sqrt(2762) = 53
"000110101",  -- sqrt(2763) = 53
"000110101",  -- sqrt(2764) = 53
"000110101",  -- sqrt(2765) = 53
"000110101",  -- sqrt(2766) = 53
"000110101",  -- sqrt(2767) = 53
"000110101",  -- sqrt(2768) = 53
"000110101",  -- sqrt(2769) = 53
"000110101",  -- sqrt(2770) = 53
"000110101",  -- sqrt(2771) = 53
"000110101",  -- sqrt(2772) = 53
"000110101",  -- sqrt(2773) = 53
"000110101",  -- sqrt(2774) = 53
"000110101",  -- sqrt(2775) = 53
"000110101",  -- sqrt(2776) = 53
"000110101",  -- sqrt(2777) = 53
"000110101",  -- sqrt(2778) = 53
"000110101",  -- sqrt(2779) = 53
"000110101",  -- sqrt(2780) = 53
"000110101",  -- sqrt(2781) = 53
"000110101",  -- sqrt(2782) = 53
"000110101",  -- sqrt(2783) = 53
"000110101",  -- sqrt(2784) = 53
"000110101",  -- sqrt(2785) = 53
"000110101",  -- sqrt(2786) = 53
"000110101",  -- sqrt(2787) = 53
"000110101",  -- sqrt(2788) = 53
"000110101",  -- sqrt(2789) = 53
"000110101",  -- sqrt(2790) = 53
"000110101",  -- sqrt(2791) = 53
"000110101",  -- sqrt(2792) = 53
"000110101",  -- sqrt(2793) = 53
"000110101",  -- sqrt(2794) = 53
"000110101",  -- sqrt(2795) = 53
"000110101",  -- sqrt(2796) = 53
"000110101",  -- sqrt(2797) = 53
"000110101",  -- sqrt(2798) = 53
"000110101",  -- sqrt(2799) = 53
"000110101",  -- sqrt(2800) = 53
"000110101",  -- sqrt(2801) = 53
"000110101",  -- sqrt(2802) = 53
"000110101",  -- sqrt(2803) = 53
"000110101",  -- sqrt(2804) = 53
"000110101",  -- sqrt(2805) = 53
"000110101",  -- sqrt(2806) = 53
"000110101",  -- sqrt(2807) = 53
"000110101",  -- sqrt(2808) = 53
"000110101",  -- sqrt(2809) = 53
"000110101",  -- sqrt(2810) = 53
"000110101",  -- sqrt(2811) = 53
"000110101",  -- sqrt(2812) = 53
"000110101",  -- sqrt(2813) = 53
"000110101",  -- sqrt(2814) = 53
"000110101",  -- sqrt(2815) = 53
"000110101",  -- sqrt(2816) = 53
"000110101",  -- sqrt(2817) = 53
"000110101",  -- sqrt(2818) = 53
"000110101",  -- sqrt(2819) = 53
"000110101",  -- sqrt(2820) = 53
"000110101",  -- sqrt(2821) = 53
"000110101",  -- sqrt(2822) = 53
"000110101",  -- sqrt(2823) = 53
"000110101",  -- sqrt(2824) = 53
"000110101",  -- sqrt(2825) = 53
"000110101",  -- sqrt(2826) = 53
"000110101",  -- sqrt(2827) = 53
"000110101",  -- sqrt(2828) = 53
"000110101",  -- sqrt(2829) = 53
"000110101",  -- sqrt(2830) = 53
"000110101",  -- sqrt(2831) = 53
"000110101",  -- sqrt(2832) = 53
"000110101",  -- sqrt(2833) = 53
"000110101",  -- sqrt(2834) = 53
"000110101",  -- sqrt(2835) = 53
"000110101",  -- sqrt(2836) = 53
"000110101",  -- sqrt(2837) = 53
"000110101",  -- sqrt(2838) = 53
"000110101",  -- sqrt(2839) = 53
"000110101",  -- sqrt(2840) = 53
"000110101",  -- sqrt(2841) = 53
"000110101",  -- sqrt(2842) = 53
"000110101",  -- sqrt(2843) = 53
"000110101",  -- sqrt(2844) = 53
"000110101",  -- sqrt(2845) = 53
"000110101",  -- sqrt(2846) = 53
"000110101",  -- sqrt(2847) = 53
"000110101",  -- sqrt(2848) = 53
"000110101",  -- sqrt(2849) = 53
"000110101",  -- sqrt(2850) = 53
"000110101",  -- sqrt(2851) = 53
"000110101",  -- sqrt(2852) = 53
"000110101",  -- sqrt(2853) = 53
"000110101",  -- sqrt(2854) = 53
"000110101",  -- sqrt(2855) = 53
"000110101",  -- sqrt(2856) = 53
"000110101",  -- sqrt(2857) = 53
"000110101",  -- sqrt(2858) = 53
"000110101",  -- sqrt(2859) = 53
"000110101",  -- sqrt(2860) = 53
"000110101",  -- sqrt(2861) = 53
"000110101",  -- sqrt(2862) = 53
"000110110",  -- sqrt(2863) = 54
"000110110",  -- sqrt(2864) = 54
"000110110",  -- sqrt(2865) = 54
"000110110",  -- sqrt(2866) = 54
"000110110",  -- sqrt(2867) = 54
"000110110",  -- sqrt(2868) = 54
"000110110",  -- sqrt(2869) = 54
"000110110",  -- sqrt(2870) = 54
"000110110",  -- sqrt(2871) = 54
"000110110",  -- sqrt(2872) = 54
"000110110",  -- sqrt(2873) = 54
"000110110",  -- sqrt(2874) = 54
"000110110",  -- sqrt(2875) = 54
"000110110",  -- sqrt(2876) = 54
"000110110",  -- sqrt(2877) = 54
"000110110",  -- sqrt(2878) = 54
"000110110",  -- sqrt(2879) = 54
"000110110",  -- sqrt(2880) = 54
"000110110",  -- sqrt(2881) = 54
"000110110",  -- sqrt(2882) = 54
"000110110",  -- sqrt(2883) = 54
"000110110",  -- sqrt(2884) = 54
"000110110",  -- sqrt(2885) = 54
"000110110",  -- sqrt(2886) = 54
"000110110",  -- sqrt(2887) = 54
"000110110",  -- sqrt(2888) = 54
"000110110",  -- sqrt(2889) = 54
"000110110",  -- sqrt(2890) = 54
"000110110",  -- sqrt(2891) = 54
"000110110",  -- sqrt(2892) = 54
"000110110",  -- sqrt(2893) = 54
"000110110",  -- sqrt(2894) = 54
"000110110",  -- sqrt(2895) = 54
"000110110",  -- sqrt(2896) = 54
"000110110",  -- sqrt(2897) = 54
"000110110",  -- sqrt(2898) = 54
"000110110",  -- sqrt(2899) = 54
"000110110",  -- sqrt(2900) = 54
"000110110",  -- sqrt(2901) = 54
"000110110",  -- sqrt(2902) = 54
"000110110",  -- sqrt(2903) = 54
"000110110",  -- sqrt(2904) = 54
"000110110",  -- sqrt(2905) = 54
"000110110",  -- sqrt(2906) = 54
"000110110",  -- sqrt(2907) = 54
"000110110",  -- sqrt(2908) = 54
"000110110",  -- sqrt(2909) = 54
"000110110",  -- sqrt(2910) = 54
"000110110",  -- sqrt(2911) = 54
"000110110",  -- sqrt(2912) = 54
"000110110",  -- sqrt(2913) = 54
"000110110",  -- sqrt(2914) = 54
"000110110",  -- sqrt(2915) = 54
"000110110",  -- sqrt(2916) = 54
"000110110",  -- sqrt(2917) = 54
"000110110",  -- sqrt(2918) = 54
"000110110",  -- sqrt(2919) = 54
"000110110",  -- sqrt(2920) = 54
"000110110",  -- sqrt(2921) = 54
"000110110",  -- sqrt(2922) = 54
"000110110",  -- sqrt(2923) = 54
"000110110",  -- sqrt(2924) = 54
"000110110",  -- sqrt(2925) = 54
"000110110",  -- sqrt(2926) = 54
"000110110",  -- sqrt(2927) = 54
"000110110",  -- sqrt(2928) = 54
"000110110",  -- sqrt(2929) = 54
"000110110",  -- sqrt(2930) = 54
"000110110",  -- sqrt(2931) = 54
"000110110",  -- sqrt(2932) = 54
"000110110",  -- sqrt(2933) = 54
"000110110",  -- sqrt(2934) = 54
"000110110",  -- sqrt(2935) = 54
"000110110",  -- sqrt(2936) = 54
"000110110",  -- sqrt(2937) = 54
"000110110",  -- sqrt(2938) = 54
"000110110",  -- sqrt(2939) = 54
"000110110",  -- sqrt(2940) = 54
"000110110",  -- sqrt(2941) = 54
"000110110",  -- sqrt(2942) = 54
"000110110",  -- sqrt(2943) = 54
"000110110",  -- sqrt(2944) = 54
"000110110",  -- sqrt(2945) = 54
"000110110",  -- sqrt(2946) = 54
"000110110",  -- sqrt(2947) = 54
"000110110",  -- sqrt(2948) = 54
"000110110",  -- sqrt(2949) = 54
"000110110",  -- sqrt(2950) = 54
"000110110",  -- sqrt(2951) = 54
"000110110",  -- sqrt(2952) = 54
"000110110",  -- sqrt(2953) = 54
"000110110",  -- sqrt(2954) = 54
"000110110",  -- sqrt(2955) = 54
"000110110",  -- sqrt(2956) = 54
"000110110",  -- sqrt(2957) = 54
"000110110",  -- sqrt(2958) = 54
"000110110",  -- sqrt(2959) = 54
"000110110",  -- sqrt(2960) = 54
"000110110",  -- sqrt(2961) = 54
"000110110",  -- sqrt(2962) = 54
"000110110",  -- sqrt(2963) = 54
"000110110",  -- sqrt(2964) = 54
"000110110",  -- sqrt(2965) = 54
"000110110",  -- sqrt(2966) = 54
"000110110",  -- sqrt(2967) = 54
"000110110",  -- sqrt(2968) = 54
"000110110",  -- sqrt(2969) = 54
"000110110",  -- sqrt(2970) = 54
"000110111",  -- sqrt(2971) = 55
"000110111",  -- sqrt(2972) = 55
"000110111",  -- sqrt(2973) = 55
"000110111",  -- sqrt(2974) = 55
"000110111",  -- sqrt(2975) = 55
"000110111",  -- sqrt(2976) = 55
"000110111",  -- sqrt(2977) = 55
"000110111",  -- sqrt(2978) = 55
"000110111",  -- sqrt(2979) = 55
"000110111",  -- sqrt(2980) = 55
"000110111",  -- sqrt(2981) = 55
"000110111",  -- sqrt(2982) = 55
"000110111",  -- sqrt(2983) = 55
"000110111",  -- sqrt(2984) = 55
"000110111",  -- sqrt(2985) = 55
"000110111",  -- sqrt(2986) = 55
"000110111",  -- sqrt(2987) = 55
"000110111",  -- sqrt(2988) = 55
"000110111",  -- sqrt(2989) = 55
"000110111",  -- sqrt(2990) = 55
"000110111",  -- sqrt(2991) = 55
"000110111",  -- sqrt(2992) = 55
"000110111",  -- sqrt(2993) = 55
"000110111",  -- sqrt(2994) = 55
"000110111",  -- sqrt(2995) = 55
"000110111",  -- sqrt(2996) = 55
"000110111",  -- sqrt(2997) = 55
"000110111",  -- sqrt(2998) = 55
"000110111",  -- sqrt(2999) = 55
"000110111",  -- sqrt(3000) = 55
"000110111",  -- sqrt(3001) = 55
"000110111",  -- sqrt(3002) = 55
"000110111",  -- sqrt(3003) = 55
"000110111",  -- sqrt(3004) = 55
"000110111",  -- sqrt(3005) = 55
"000110111",  -- sqrt(3006) = 55
"000110111",  -- sqrt(3007) = 55
"000110111",  -- sqrt(3008) = 55
"000110111",  -- sqrt(3009) = 55
"000110111",  -- sqrt(3010) = 55
"000110111",  -- sqrt(3011) = 55
"000110111",  -- sqrt(3012) = 55
"000110111",  -- sqrt(3013) = 55
"000110111",  -- sqrt(3014) = 55
"000110111",  -- sqrt(3015) = 55
"000110111",  -- sqrt(3016) = 55
"000110111",  -- sqrt(3017) = 55
"000110111",  -- sqrt(3018) = 55
"000110111",  -- sqrt(3019) = 55
"000110111",  -- sqrt(3020) = 55
"000110111",  -- sqrt(3021) = 55
"000110111",  -- sqrt(3022) = 55
"000110111",  -- sqrt(3023) = 55
"000110111",  -- sqrt(3024) = 55
"000110111",  -- sqrt(3025) = 55
"000110111",  -- sqrt(3026) = 55
"000110111",  -- sqrt(3027) = 55
"000110111",  -- sqrt(3028) = 55
"000110111",  -- sqrt(3029) = 55
"000110111",  -- sqrt(3030) = 55
"000110111",  -- sqrt(3031) = 55
"000110111",  -- sqrt(3032) = 55
"000110111",  -- sqrt(3033) = 55
"000110111",  -- sqrt(3034) = 55
"000110111",  -- sqrt(3035) = 55
"000110111",  -- sqrt(3036) = 55
"000110111",  -- sqrt(3037) = 55
"000110111",  -- sqrt(3038) = 55
"000110111",  -- sqrt(3039) = 55
"000110111",  -- sqrt(3040) = 55
"000110111",  -- sqrt(3041) = 55
"000110111",  -- sqrt(3042) = 55
"000110111",  -- sqrt(3043) = 55
"000110111",  -- sqrt(3044) = 55
"000110111",  -- sqrt(3045) = 55
"000110111",  -- sqrt(3046) = 55
"000110111",  -- sqrt(3047) = 55
"000110111",  -- sqrt(3048) = 55
"000110111",  -- sqrt(3049) = 55
"000110111",  -- sqrt(3050) = 55
"000110111",  -- sqrt(3051) = 55
"000110111",  -- sqrt(3052) = 55
"000110111",  -- sqrt(3053) = 55
"000110111",  -- sqrt(3054) = 55
"000110111",  -- sqrt(3055) = 55
"000110111",  -- sqrt(3056) = 55
"000110111",  -- sqrt(3057) = 55
"000110111",  -- sqrt(3058) = 55
"000110111",  -- sqrt(3059) = 55
"000110111",  -- sqrt(3060) = 55
"000110111",  -- sqrt(3061) = 55
"000110111",  -- sqrt(3062) = 55
"000110111",  -- sqrt(3063) = 55
"000110111",  -- sqrt(3064) = 55
"000110111",  -- sqrt(3065) = 55
"000110111",  -- sqrt(3066) = 55
"000110111",  -- sqrt(3067) = 55
"000110111",  -- sqrt(3068) = 55
"000110111",  -- sqrt(3069) = 55
"000110111",  -- sqrt(3070) = 55
"000110111",  -- sqrt(3071) = 55
"000110111",  -- sqrt(3072) = 55
"000110111",  -- sqrt(3073) = 55
"000110111",  -- sqrt(3074) = 55
"000110111",  -- sqrt(3075) = 55
"000110111",  -- sqrt(3076) = 55
"000110111",  -- sqrt(3077) = 55
"000110111",  -- sqrt(3078) = 55
"000110111",  -- sqrt(3079) = 55
"000110111",  -- sqrt(3080) = 55
"000111000",  -- sqrt(3081) = 56
"000111000",  -- sqrt(3082) = 56
"000111000",  -- sqrt(3083) = 56
"000111000",  -- sqrt(3084) = 56
"000111000",  -- sqrt(3085) = 56
"000111000",  -- sqrt(3086) = 56
"000111000",  -- sqrt(3087) = 56
"000111000",  -- sqrt(3088) = 56
"000111000",  -- sqrt(3089) = 56
"000111000",  -- sqrt(3090) = 56
"000111000",  -- sqrt(3091) = 56
"000111000",  -- sqrt(3092) = 56
"000111000",  -- sqrt(3093) = 56
"000111000",  -- sqrt(3094) = 56
"000111000",  -- sqrt(3095) = 56
"000111000",  -- sqrt(3096) = 56
"000111000",  -- sqrt(3097) = 56
"000111000",  -- sqrt(3098) = 56
"000111000",  -- sqrt(3099) = 56
"000111000",  -- sqrt(3100) = 56
"000111000",  -- sqrt(3101) = 56
"000111000",  -- sqrt(3102) = 56
"000111000",  -- sqrt(3103) = 56
"000111000",  -- sqrt(3104) = 56
"000111000",  -- sqrt(3105) = 56
"000111000",  -- sqrt(3106) = 56
"000111000",  -- sqrt(3107) = 56
"000111000",  -- sqrt(3108) = 56
"000111000",  -- sqrt(3109) = 56
"000111000",  -- sqrt(3110) = 56
"000111000",  -- sqrt(3111) = 56
"000111000",  -- sqrt(3112) = 56
"000111000",  -- sqrt(3113) = 56
"000111000",  -- sqrt(3114) = 56
"000111000",  -- sqrt(3115) = 56
"000111000",  -- sqrt(3116) = 56
"000111000",  -- sqrt(3117) = 56
"000111000",  -- sqrt(3118) = 56
"000111000",  -- sqrt(3119) = 56
"000111000",  -- sqrt(3120) = 56
"000111000",  -- sqrt(3121) = 56
"000111000",  -- sqrt(3122) = 56
"000111000",  -- sqrt(3123) = 56
"000111000",  -- sqrt(3124) = 56
"000111000",  -- sqrt(3125) = 56
"000111000",  -- sqrt(3126) = 56
"000111000",  -- sqrt(3127) = 56
"000111000",  -- sqrt(3128) = 56
"000111000",  -- sqrt(3129) = 56
"000111000",  -- sqrt(3130) = 56
"000111000",  -- sqrt(3131) = 56
"000111000",  -- sqrt(3132) = 56
"000111000",  -- sqrt(3133) = 56
"000111000",  -- sqrt(3134) = 56
"000111000",  -- sqrt(3135) = 56
"000111000",  -- sqrt(3136) = 56
"000111000",  -- sqrt(3137) = 56
"000111000",  -- sqrt(3138) = 56
"000111000",  -- sqrt(3139) = 56
"000111000",  -- sqrt(3140) = 56
"000111000",  -- sqrt(3141) = 56
"000111000",  -- sqrt(3142) = 56
"000111000",  -- sqrt(3143) = 56
"000111000",  -- sqrt(3144) = 56
"000111000",  -- sqrt(3145) = 56
"000111000",  -- sqrt(3146) = 56
"000111000",  -- sqrt(3147) = 56
"000111000",  -- sqrt(3148) = 56
"000111000",  -- sqrt(3149) = 56
"000111000",  -- sqrt(3150) = 56
"000111000",  -- sqrt(3151) = 56
"000111000",  -- sqrt(3152) = 56
"000111000",  -- sqrt(3153) = 56
"000111000",  -- sqrt(3154) = 56
"000111000",  -- sqrt(3155) = 56
"000111000",  -- sqrt(3156) = 56
"000111000",  -- sqrt(3157) = 56
"000111000",  -- sqrt(3158) = 56
"000111000",  -- sqrt(3159) = 56
"000111000",  -- sqrt(3160) = 56
"000111000",  -- sqrt(3161) = 56
"000111000",  -- sqrt(3162) = 56
"000111000",  -- sqrt(3163) = 56
"000111000",  -- sqrt(3164) = 56
"000111000",  -- sqrt(3165) = 56
"000111000",  -- sqrt(3166) = 56
"000111000",  -- sqrt(3167) = 56
"000111000",  -- sqrt(3168) = 56
"000111000",  -- sqrt(3169) = 56
"000111000",  -- sqrt(3170) = 56
"000111000",  -- sqrt(3171) = 56
"000111000",  -- sqrt(3172) = 56
"000111000",  -- sqrt(3173) = 56
"000111000",  -- sqrt(3174) = 56
"000111000",  -- sqrt(3175) = 56
"000111000",  -- sqrt(3176) = 56
"000111000",  -- sqrt(3177) = 56
"000111000",  -- sqrt(3178) = 56
"000111000",  -- sqrt(3179) = 56
"000111000",  -- sqrt(3180) = 56
"000111000",  -- sqrt(3181) = 56
"000111000",  -- sqrt(3182) = 56
"000111000",  -- sqrt(3183) = 56
"000111000",  -- sqrt(3184) = 56
"000111000",  -- sqrt(3185) = 56
"000111000",  -- sqrt(3186) = 56
"000111000",  -- sqrt(3187) = 56
"000111000",  -- sqrt(3188) = 56
"000111000",  -- sqrt(3189) = 56
"000111000",  -- sqrt(3190) = 56
"000111000",  -- sqrt(3191) = 56
"000111000",  -- sqrt(3192) = 56
"000111001",  -- sqrt(3193) = 57
"000111001",  -- sqrt(3194) = 57
"000111001",  -- sqrt(3195) = 57
"000111001",  -- sqrt(3196) = 57
"000111001",  -- sqrt(3197) = 57
"000111001",  -- sqrt(3198) = 57
"000111001",  -- sqrt(3199) = 57
"000111001",  -- sqrt(3200) = 57
"000111001",  -- sqrt(3201) = 57
"000111001",  -- sqrt(3202) = 57
"000111001",  -- sqrt(3203) = 57
"000111001",  -- sqrt(3204) = 57
"000111001",  -- sqrt(3205) = 57
"000111001",  -- sqrt(3206) = 57
"000111001",  -- sqrt(3207) = 57
"000111001",  -- sqrt(3208) = 57
"000111001",  -- sqrt(3209) = 57
"000111001",  -- sqrt(3210) = 57
"000111001",  -- sqrt(3211) = 57
"000111001",  -- sqrt(3212) = 57
"000111001",  -- sqrt(3213) = 57
"000111001",  -- sqrt(3214) = 57
"000111001",  -- sqrt(3215) = 57
"000111001",  -- sqrt(3216) = 57
"000111001",  -- sqrt(3217) = 57
"000111001",  -- sqrt(3218) = 57
"000111001",  -- sqrt(3219) = 57
"000111001",  -- sqrt(3220) = 57
"000111001",  -- sqrt(3221) = 57
"000111001",  -- sqrt(3222) = 57
"000111001",  -- sqrt(3223) = 57
"000111001",  -- sqrt(3224) = 57
"000111001",  -- sqrt(3225) = 57
"000111001",  -- sqrt(3226) = 57
"000111001",  -- sqrt(3227) = 57
"000111001",  -- sqrt(3228) = 57
"000111001",  -- sqrt(3229) = 57
"000111001",  -- sqrt(3230) = 57
"000111001",  -- sqrt(3231) = 57
"000111001",  -- sqrt(3232) = 57
"000111001",  -- sqrt(3233) = 57
"000111001",  -- sqrt(3234) = 57
"000111001",  -- sqrt(3235) = 57
"000111001",  -- sqrt(3236) = 57
"000111001",  -- sqrt(3237) = 57
"000111001",  -- sqrt(3238) = 57
"000111001",  -- sqrt(3239) = 57
"000111001",  -- sqrt(3240) = 57
"000111001",  -- sqrt(3241) = 57
"000111001",  -- sqrt(3242) = 57
"000111001",  -- sqrt(3243) = 57
"000111001",  -- sqrt(3244) = 57
"000111001",  -- sqrt(3245) = 57
"000111001",  -- sqrt(3246) = 57
"000111001",  -- sqrt(3247) = 57
"000111001",  -- sqrt(3248) = 57
"000111001",  -- sqrt(3249) = 57
"000111001",  -- sqrt(3250) = 57
"000111001",  -- sqrt(3251) = 57
"000111001",  -- sqrt(3252) = 57
"000111001",  -- sqrt(3253) = 57
"000111001",  -- sqrt(3254) = 57
"000111001",  -- sqrt(3255) = 57
"000111001",  -- sqrt(3256) = 57
"000111001",  -- sqrt(3257) = 57
"000111001",  -- sqrt(3258) = 57
"000111001",  -- sqrt(3259) = 57
"000111001",  -- sqrt(3260) = 57
"000111001",  -- sqrt(3261) = 57
"000111001",  -- sqrt(3262) = 57
"000111001",  -- sqrt(3263) = 57
"000111001",  -- sqrt(3264) = 57
"000111001",  -- sqrt(3265) = 57
"000111001",  -- sqrt(3266) = 57
"000111001",  -- sqrt(3267) = 57
"000111001",  -- sqrt(3268) = 57
"000111001",  -- sqrt(3269) = 57
"000111001",  -- sqrt(3270) = 57
"000111001",  -- sqrt(3271) = 57
"000111001",  -- sqrt(3272) = 57
"000111001",  -- sqrt(3273) = 57
"000111001",  -- sqrt(3274) = 57
"000111001",  -- sqrt(3275) = 57
"000111001",  -- sqrt(3276) = 57
"000111001",  -- sqrt(3277) = 57
"000111001",  -- sqrt(3278) = 57
"000111001",  -- sqrt(3279) = 57
"000111001",  -- sqrt(3280) = 57
"000111001",  -- sqrt(3281) = 57
"000111001",  -- sqrt(3282) = 57
"000111001",  -- sqrt(3283) = 57
"000111001",  -- sqrt(3284) = 57
"000111001",  -- sqrt(3285) = 57
"000111001",  -- sqrt(3286) = 57
"000111001",  -- sqrt(3287) = 57
"000111001",  -- sqrt(3288) = 57
"000111001",  -- sqrt(3289) = 57
"000111001",  -- sqrt(3290) = 57
"000111001",  -- sqrt(3291) = 57
"000111001",  -- sqrt(3292) = 57
"000111001",  -- sqrt(3293) = 57
"000111001",  -- sqrt(3294) = 57
"000111001",  -- sqrt(3295) = 57
"000111001",  -- sqrt(3296) = 57
"000111001",  -- sqrt(3297) = 57
"000111001",  -- sqrt(3298) = 57
"000111001",  -- sqrt(3299) = 57
"000111001",  -- sqrt(3300) = 57
"000111001",  -- sqrt(3301) = 57
"000111001",  -- sqrt(3302) = 57
"000111001",  -- sqrt(3303) = 57
"000111001",  -- sqrt(3304) = 57
"000111001",  -- sqrt(3305) = 57
"000111001",  -- sqrt(3306) = 57
"000111010",  -- sqrt(3307) = 58
"000111010",  -- sqrt(3308) = 58
"000111010",  -- sqrt(3309) = 58
"000111010",  -- sqrt(3310) = 58
"000111010",  -- sqrt(3311) = 58
"000111010",  -- sqrt(3312) = 58
"000111010",  -- sqrt(3313) = 58
"000111010",  -- sqrt(3314) = 58
"000111010",  -- sqrt(3315) = 58
"000111010",  -- sqrt(3316) = 58
"000111010",  -- sqrt(3317) = 58
"000111010",  -- sqrt(3318) = 58
"000111010",  -- sqrt(3319) = 58
"000111010",  -- sqrt(3320) = 58
"000111010",  -- sqrt(3321) = 58
"000111010",  -- sqrt(3322) = 58
"000111010",  -- sqrt(3323) = 58
"000111010",  -- sqrt(3324) = 58
"000111010",  -- sqrt(3325) = 58
"000111010",  -- sqrt(3326) = 58
"000111010",  -- sqrt(3327) = 58
"000111010",  -- sqrt(3328) = 58
"000111010",  -- sqrt(3329) = 58
"000111010",  -- sqrt(3330) = 58
"000111010",  -- sqrt(3331) = 58
"000111010",  -- sqrt(3332) = 58
"000111010",  -- sqrt(3333) = 58
"000111010",  -- sqrt(3334) = 58
"000111010",  -- sqrt(3335) = 58
"000111010",  -- sqrt(3336) = 58
"000111010",  -- sqrt(3337) = 58
"000111010",  -- sqrt(3338) = 58
"000111010",  -- sqrt(3339) = 58
"000111010",  -- sqrt(3340) = 58
"000111010",  -- sqrt(3341) = 58
"000111010",  -- sqrt(3342) = 58
"000111010",  -- sqrt(3343) = 58
"000111010",  -- sqrt(3344) = 58
"000111010",  -- sqrt(3345) = 58
"000111010",  -- sqrt(3346) = 58
"000111010",  -- sqrt(3347) = 58
"000111010",  -- sqrt(3348) = 58
"000111010",  -- sqrt(3349) = 58
"000111010",  -- sqrt(3350) = 58
"000111010",  -- sqrt(3351) = 58
"000111010",  -- sqrt(3352) = 58
"000111010",  -- sqrt(3353) = 58
"000111010",  -- sqrt(3354) = 58
"000111010",  -- sqrt(3355) = 58
"000111010",  -- sqrt(3356) = 58
"000111010",  -- sqrt(3357) = 58
"000111010",  -- sqrt(3358) = 58
"000111010",  -- sqrt(3359) = 58
"000111010",  -- sqrt(3360) = 58
"000111010",  -- sqrt(3361) = 58
"000111010",  -- sqrt(3362) = 58
"000111010",  -- sqrt(3363) = 58
"000111010",  -- sqrt(3364) = 58
"000111010",  -- sqrt(3365) = 58
"000111010",  -- sqrt(3366) = 58
"000111010",  -- sqrt(3367) = 58
"000111010",  -- sqrt(3368) = 58
"000111010",  -- sqrt(3369) = 58
"000111010",  -- sqrt(3370) = 58
"000111010",  -- sqrt(3371) = 58
"000111010",  -- sqrt(3372) = 58
"000111010",  -- sqrt(3373) = 58
"000111010",  -- sqrt(3374) = 58
"000111010",  -- sqrt(3375) = 58
"000111010",  -- sqrt(3376) = 58
"000111010",  -- sqrt(3377) = 58
"000111010",  -- sqrt(3378) = 58
"000111010",  -- sqrt(3379) = 58
"000111010",  -- sqrt(3380) = 58
"000111010",  -- sqrt(3381) = 58
"000111010",  -- sqrt(3382) = 58
"000111010",  -- sqrt(3383) = 58
"000111010",  -- sqrt(3384) = 58
"000111010",  -- sqrt(3385) = 58
"000111010",  -- sqrt(3386) = 58
"000111010",  -- sqrt(3387) = 58
"000111010",  -- sqrt(3388) = 58
"000111010",  -- sqrt(3389) = 58
"000111010",  -- sqrt(3390) = 58
"000111010",  -- sqrt(3391) = 58
"000111010",  -- sqrt(3392) = 58
"000111010",  -- sqrt(3393) = 58
"000111010",  -- sqrt(3394) = 58
"000111010",  -- sqrt(3395) = 58
"000111010",  -- sqrt(3396) = 58
"000111010",  -- sqrt(3397) = 58
"000111010",  -- sqrt(3398) = 58
"000111010",  -- sqrt(3399) = 58
"000111010",  -- sqrt(3400) = 58
"000111010",  -- sqrt(3401) = 58
"000111010",  -- sqrt(3402) = 58
"000111010",  -- sqrt(3403) = 58
"000111010",  -- sqrt(3404) = 58
"000111010",  -- sqrt(3405) = 58
"000111010",  -- sqrt(3406) = 58
"000111010",  -- sqrt(3407) = 58
"000111010",  -- sqrt(3408) = 58
"000111010",  -- sqrt(3409) = 58
"000111010",  -- sqrt(3410) = 58
"000111010",  -- sqrt(3411) = 58
"000111010",  -- sqrt(3412) = 58
"000111010",  -- sqrt(3413) = 58
"000111010",  -- sqrt(3414) = 58
"000111010",  -- sqrt(3415) = 58
"000111010",  -- sqrt(3416) = 58
"000111010",  -- sqrt(3417) = 58
"000111010",  -- sqrt(3418) = 58
"000111010",  -- sqrt(3419) = 58
"000111010",  -- sqrt(3420) = 58
"000111010",  -- sqrt(3421) = 58
"000111010",  -- sqrt(3422) = 58
"000111011",  -- sqrt(3423) = 59
"000111011",  -- sqrt(3424) = 59
"000111011",  -- sqrt(3425) = 59
"000111011",  -- sqrt(3426) = 59
"000111011",  -- sqrt(3427) = 59
"000111011",  -- sqrt(3428) = 59
"000111011",  -- sqrt(3429) = 59
"000111011",  -- sqrt(3430) = 59
"000111011",  -- sqrt(3431) = 59
"000111011",  -- sqrt(3432) = 59
"000111011",  -- sqrt(3433) = 59
"000111011",  -- sqrt(3434) = 59
"000111011",  -- sqrt(3435) = 59
"000111011",  -- sqrt(3436) = 59
"000111011",  -- sqrt(3437) = 59
"000111011",  -- sqrt(3438) = 59
"000111011",  -- sqrt(3439) = 59
"000111011",  -- sqrt(3440) = 59
"000111011",  -- sqrt(3441) = 59
"000111011",  -- sqrt(3442) = 59
"000111011",  -- sqrt(3443) = 59
"000111011",  -- sqrt(3444) = 59
"000111011",  -- sqrt(3445) = 59
"000111011",  -- sqrt(3446) = 59
"000111011",  -- sqrt(3447) = 59
"000111011",  -- sqrt(3448) = 59
"000111011",  -- sqrt(3449) = 59
"000111011",  -- sqrt(3450) = 59
"000111011",  -- sqrt(3451) = 59
"000111011",  -- sqrt(3452) = 59
"000111011",  -- sqrt(3453) = 59
"000111011",  -- sqrt(3454) = 59
"000111011",  -- sqrt(3455) = 59
"000111011",  -- sqrt(3456) = 59
"000111011",  -- sqrt(3457) = 59
"000111011",  -- sqrt(3458) = 59
"000111011",  -- sqrt(3459) = 59
"000111011",  -- sqrt(3460) = 59
"000111011",  -- sqrt(3461) = 59
"000111011",  -- sqrt(3462) = 59
"000111011",  -- sqrt(3463) = 59
"000111011",  -- sqrt(3464) = 59
"000111011",  -- sqrt(3465) = 59
"000111011",  -- sqrt(3466) = 59
"000111011",  -- sqrt(3467) = 59
"000111011",  -- sqrt(3468) = 59
"000111011",  -- sqrt(3469) = 59
"000111011",  -- sqrt(3470) = 59
"000111011",  -- sqrt(3471) = 59
"000111011",  -- sqrt(3472) = 59
"000111011",  -- sqrt(3473) = 59
"000111011",  -- sqrt(3474) = 59
"000111011",  -- sqrt(3475) = 59
"000111011",  -- sqrt(3476) = 59
"000111011",  -- sqrt(3477) = 59
"000111011",  -- sqrt(3478) = 59
"000111011",  -- sqrt(3479) = 59
"000111011",  -- sqrt(3480) = 59
"000111011",  -- sqrt(3481) = 59
"000111011",  -- sqrt(3482) = 59
"000111011",  -- sqrt(3483) = 59
"000111011",  -- sqrt(3484) = 59
"000111011",  -- sqrt(3485) = 59
"000111011",  -- sqrt(3486) = 59
"000111011",  -- sqrt(3487) = 59
"000111011",  -- sqrt(3488) = 59
"000111011",  -- sqrt(3489) = 59
"000111011",  -- sqrt(3490) = 59
"000111011",  -- sqrt(3491) = 59
"000111011",  -- sqrt(3492) = 59
"000111011",  -- sqrt(3493) = 59
"000111011",  -- sqrt(3494) = 59
"000111011",  -- sqrt(3495) = 59
"000111011",  -- sqrt(3496) = 59
"000111011",  -- sqrt(3497) = 59
"000111011",  -- sqrt(3498) = 59
"000111011",  -- sqrt(3499) = 59
"000111011",  -- sqrt(3500) = 59
"000111011",  -- sqrt(3501) = 59
"000111011",  -- sqrt(3502) = 59
"000111011",  -- sqrt(3503) = 59
"000111011",  -- sqrt(3504) = 59
"000111011",  -- sqrt(3505) = 59
"000111011",  -- sqrt(3506) = 59
"000111011",  -- sqrt(3507) = 59
"000111011",  -- sqrt(3508) = 59
"000111011",  -- sqrt(3509) = 59
"000111011",  -- sqrt(3510) = 59
"000111011",  -- sqrt(3511) = 59
"000111011",  -- sqrt(3512) = 59
"000111011",  -- sqrt(3513) = 59
"000111011",  -- sqrt(3514) = 59
"000111011",  -- sqrt(3515) = 59
"000111011",  -- sqrt(3516) = 59
"000111011",  -- sqrt(3517) = 59
"000111011",  -- sqrt(3518) = 59
"000111011",  -- sqrt(3519) = 59
"000111011",  -- sqrt(3520) = 59
"000111011",  -- sqrt(3521) = 59
"000111011",  -- sqrt(3522) = 59
"000111011",  -- sqrt(3523) = 59
"000111011",  -- sqrt(3524) = 59
"000111011",  -- sqrt(3525) = 59
"000111011",  -- sqrt(3526) = 59
"000111011",  -- sqrt(3527) = 59
"000111011",  -- sqrt(3528) = 59
"000111011",  -- sqrt(3529) = 59
"000111011",  -- sqrt(3530) = 59
"000111011",  -- sqrt(3531) = 59
"000111011",  -- sqrt(3532) = 59
"000111011",  -- sqrt(3533) = 59
"000111011",  -- sqrt(3534) = 59
"000111011",  -- sqrt(3535) = 59
"000111011",  -- sqrt(3536) = 59
"000111011",  -- sqrt(3537) = 59
"000111011",  -- sqrt(3538) = 59
"000111011",  -- sqrt(3539) = 59
"000111011",  -- sqrt(3540) = 59
"000111100",  -- sqrt(3541) = 60
"000111100",  -- sqrt(3542) = 60
"000111100",  -- sqrt(3543) = 60
"000111100",  -- sqrt(3544) = 60
"000111100",  -- sqrt(3545) = 60
"000111100",  -- sqrt(3546) = 60
"000111100",  -- sqrt(3547) = 60
"000111100",  -- sqrt(3548) = 60
"000111100",  -- sqrt(3549) = 60
"000111100",  -- sqrt(3550) = 60
"000111100",  -- sqrt(3551) = 60
"000111100",  -- sqrt(3552) = 60
"000111100",  -- sqrt(3553) = 60
"000111100",  -- sqrt(3554) = 60
"000111100",  -- sqrt(3555) = 60
"000111100",  -- sqrt(3556) = 60
"000111100",  -- sqrt(3557) = 60
"000111100",  -- sqrt(3558) = 60
"000111100",  -- sqrt(3559) = 60
"000111100",  -- sqrt(3560) = 60
"000111100",  -- sqrt(3561) = 60
"000111100",  -- sqrt(3562) = 60
"000111100",  -- sqrt(3563) = 60
"000111100",  -- sqrt(3564) = 60
"000111100",  -- sqrt(3565) = 60
"000111100",  -- sqrt(3566) = 60
"000111100",  -- sqrt(3567) = 60
"000111100",  -- sqrt(3568) = 60
"000111100",  -- sqrt(3569) = 60
"000111100",  -- sqrt(3570) = 60
"000111100",  -- sqrt(3571) = 60
"000111100",  -- sqrt(3572) = 60
"000111100",  -- sqrt(3573) = 60
"000111100",  -- sqrt(3574) = 60
"000111100",  -- sqrt(3575) = 60
"000111100",  -- sqrt(3576) = 60
"000111100",  -- sqrt(3577) = 60
"000111100",  -- sqrt(3578) = 60
"000111100",  -- sqrt(3579) = 60
"000111100",  -- sqrt(3580) = 60
"000111100",  -- sqrt(3581) = 60
"000111100",  -- sqrt(3582) = 60
"000111100",  -- sqrt(3583) = 60
"000111100",  -- sqrt(3584) = 60
"000111100",  -- sqrt(3585) = 60
"000111100",  -- sqrt(3586) = 60
"000111100",  -- sqrt(3587) = 60
"000111100",  -- sqrt(3588) = 60
"000111100",  -- sqrt(3589) = 60
"000111100",  -- sqrt(3590) = 60
"000111100",  -- sqrt(3591) = 60
"000111100",  -- sqrt(3592) = 60
"000111100",  -- sqrt(3593) = 60
"000111100",  -- sqrt(3594) = 60
"000111100",  -- sqrt(3595) = 60
"000111100",  -- sqrt(3596) = 60
"000111100",  -- sqrt(3597) = 60
"000111100",  -- sqrt(3598) = 60
"000111100",  -- sqrt(3599) = 60
"000111100",  -- sqrt(3600) = 60
"000111100",  -- sqrt(3601) = 60
"000111100",  -- sqrt(3602) = 60
"000111100",  -- sqrt(3603) = 60
"000111100",  -- sqrt(3604) = 60
"000111100",  -- sqrt(3605) = 60
"000111100",  -- sqrt(3606) = 60
"000111100",  -- sqrt(3607) = 60
"000111100",  -- sqrt(3608) = 60
"000111100",  -- sqrt(3609) = 60
"000111100",  -- sqrt(3610) = 60
"000111100",  -- sqrt(3611) = 60
"000111100",  -- sqrt(3612) = 60
"000111100",  -- sqrt(3613) = 60
"000111100",  -- sqrt(3614) = 60
"000111100",  -- sqrt(3615) = 60
"000111100",  -- sqrt(3616) = 60
"000111100",  -- sqrt(3617) = 60
"000111100",  -- sqrt(3618) = 60
"000111100",  -- sqrt(3619) = 60
"000111100",  -- sqrt(3620) = 60
"000111100",  -- sqrt(3621) = 60
"000111100",  -- sqrt(3622) = 60
"000111100",  -- sqrt(3623) = 60
"000111100",  -- sqrt(3624) = 60
"000111100",  -- sqrt(3625) = 60
"000111100",  -- sqrt(3626) = 60
"000111100",  -- sqrt(3627) = 60
"000111100",  -- sqrt(3628) = 60
"000111100",  -- sqrt(3629) = 60
"000111100",  -- sqrt(3630) = 60
"000111100",  -- sqrt(3631) = 60
"000111100",  -- sqrt(3632) = 60
"000111100",  -- sqrt(3633) = 60
"000111100",  -- sqrt(3634) = 60
"000111100",  -- sqrt(3635) = 60
"000111100",  -- sqrt(3636) = 60
"000111100",  -- sqrt(3637) = 60
"000111100",  -- sqrt(3638) = 60
"000111100",  -- sqrt(3639) = 60
"000111100",  -- sqrt(3640) = 60
"000111100",  -- sqrt(3641) = 60
"000111100",  -- sqrt(3642) = 60
"000111100",  -- sqrt(3643) = 60
"000111100",  -- sqrt(3644) = 60
"000111100",  -- sqrt(3645) = 60
"000111100",  -- sqrt(3646) = 60
"000111100",  -- sqrt(3647) = 60
"000111100",  -- sqrt(3648) = 60
"000111100",  -- sqrt(3649) = 60
"000111100",  -- sqrt(3650) = 60
"000111100",  -- sqrt(3651) = 60
"000111100",  -- sqrt(3652) = 60
"000111100",  -- sqrt(3653) = 60
"000111100",  -- sqrt(3654) = 60
"000111100",  -- sqrt(3655) = 60
"000111100",  -- sqrt(3656) = 60
"000111100",  -- sqrt(3657) = 60
"000111100",  -- sqrt(3658) = 60
"000111100",  -- sqrt(3659) = 60
"000111100",  -- sqrt(3660) = 60
"000111101",  -- sqrt(3661) = 61
"000111101",  -- sqrt(3662) = 61
"000111101",  -- sqrt(3663) = 61
"000111101",  -- sqrt(3664) = 61
"000111101",  -- sqrt(3665) = 61
"000111101",  -- sqrt(3666) = 61
"000111101",  -- sqrt(3667) = 61
"000111101",  -- sqrt(3668) = 61
"000111101",  -- sqrt(3669) = 61
"000111101",  -- sqrt(3670) = 61
"000111101",  -- sqrt(3671) = 61
"000111101",  -- sqrt(3672) = 61
"000111101",  -- sqrt(3673) = 61
"000111101",  -- sqrt(3674) = 61
"000111101",  -- sqrt(3675) = 61
"000111101",  -- sqrt(3676) = 61
"000111101",  -- sqrt(3677) = 61
"000111101",  -- sqrt(3678) = 61
"000111101",  -- sqrt(3679) = 61
"000111101",  -- sqrt(3680) = 61
"000111101",  -- sqrt(3681) = 61
"000111101",  -- sqrt(3682) = 61
"000111101",  -- sqrt(3683) = 61
"000111101",  -- sqrt(3684) = 61
"000111101",  -- sqrt(3685) = 61
"000111101",  -- sqrt(3686) = 61
"000111101",  -- sqrt(3687) = 61
"000111101",  -- sqrt(3688) = 61
"000111101",  -- sqrt(3689) = 61
"000111101",  -- sqrt(3690) = 61
"000111101",  -- sqrt(3691) = 61
"000111101",  -- sqrt(3692) = 61
"000111101",  -- sqrt(3693) = 61
"000111101",  -- sqrt(3694) = 61
"000111101",  -- sqrt(3695) = 61
"000111101",  -- sqrt(3696) = 61
"000111101",  -- sqrt(3697) = 61
"000111101",  -- sqrt(3698) = 61
"000111101",  -- sqrt(3699) = 61
"000111101",  -- sqrt(3700) = 61
"000111101",  -- sqrt(3701) = 61
"000111101",  -- sqrt(3702) = 61
"000111101",  -- sqrt(3703) = 61
"000111101",  -- sqrt(3704) = 61
"000111101",  -- sqrt(3705) = 61
"000111101",  -- sqrt(3706) = 61
"000111101",  -- sqrt(3707) = 61
"000111101",  -- sqrt(3708) = 61
"000111101",  -- sqrt(3709) = 61
"000111101",  -- sqrt(3710) = 61
"000111101",  -- sqrt(3711) = 61
"000111101",  -- sqrt(3712) = 61
"000111101",  -- sqrt(3713) = 61
"000111101",  -- sqrt(3714) = 61
"000111101",  -- sqrt(3715) = 61
"000111101",  -- sqrt(3716) = 61
"000111101",  -- sqrt(3717) = 61
"000111101",  -- sqrt(3718) = 61
"000111101",  -- sqrt(3719) = 61
"000111101",  -- sqrt(3720) = 61
"000111101",  -- sqrt(3721) = 61
"000111101",  -- sqrt(3722) = 61
"000111101",  -- sqrt(3723) = 61
"000111101",  -- sqrt(3724) = 61
"000111101",  -- sqrt(3725) = 61
"000111101",  -- sqrt(3726) = 61
"000111101",  -- sqrt(3727) = 61
"000111101",  -- sqrt(3728) = 61
"000111101",  -- sqrt(3729) = 61
"000111101",  -- sqrt(3730) = 61
"000111101",  -- sqrt(3731) = 61
"000111101",  -- sqrt(3732) = 61
"000111101",  -- sqrt(3733) = 61
"000111101",  -- sqrt(3734) = 61
"000111101",  -- sqrt(3735) = 61
"000111101",  -- sqrt(3736) = 61
"000111101",  -- sqrt(3737) = 61
"000111101",  -- sqrt(3738) = 61
"000111101",  -- sqrt(3739) = 61
"000111101",  -- sqrt(3740) = 61
"000111101",  -- sqrt(3741) = 61
"000111101",  -- sqrt(3742) = 61
"000111101",  -- sqrt(3743) = 61
"000111101",  -- sqrt(3744) = 61
"000111101",  -- sqrt(3745) = 61
"000111101",  -- sqrt(3746) = 61
"000111101",  -- sqrt(3747) = 61
"000111101",  -- sqrt(3748) = 61
"000111101",  -- sqrt(3749) = 61
"000111101",  -- sqrt(3750) = 61
"000111101",  -- sqrt(3751) = 61
"000111101",  -- sqrt(3752) = 61
"000111101",  -- sqrt(3753) = 61
"000111101",  -- sqrt(3754) = 61
"000111101",  -- sqrt(3755) = 61
"000111101",  -- sqrt(3756) = 61
"000111101",  -- sqrt(3757) = 61
"000111101",  -- sqrt(3758) = 61
"000111101",  -- sqrt(3759) = 61
"000111101",  -- sqrt(3760) = 61
"000111101",  -- sqrt(3761) = 61
"000111101",  -- sqrt(3762) = 61
"000111101",  -- sqrt(3763) = 61
"000111101",  -- sqrt(3764) = 61
"000111101",  -- sqrt(3765) = 61
"000111101",  -- sqrt(3766) = 61
"000111101",  -- sqrt(3767) = 61
"000111101",  -- sqrt(3768) = 61
"000111101",  -- sqrt(3769) = 61
"000111101",  -- sqrt(3770) = 61
"000111101",  -- sqrt(3771) = 61
"000111101",  -- sqrt(3772) = 61
"000111101",  -- sqrt(3773) = 61
"000111101",  -- sqrt(3774) = 61
"000111101",  -- sqrt(3775) = 61
"000111101",  -- sqrt(3776) = 61
"000111101",  -- sqrt(3777) = 61
"000111101",  -- sqrt(3778) = 61
"000111101",  -- sqrt(3779) = 61
"000111101",  -- sqrt(3780) = 61
"000111101",  -- sqrt(3781) = 61
"000111101",  -- sqrt(3782) = 61
"000111110",  -- sqrt(3783) = 62
"000111110",  -- sqrt(3784) = 62
"000111110",  -- sqrt(3785) = 62
"000111110",  -- sqrt(3786) = 62
"000111110",  -- sqrt(3787) = 62
"000111110",  -- sqrt(3788) = 62
"000111110",  -- sqrt(3789) = 62
"000111110",  -- sqrt(3790) = 62
"000111110",  -- sqrt(3791) = 62
"000111110",  -- sqrt(3792) = 62
"000111110",  -- sqrt(3793) = 62
"000111110",  -- sqrt(3794) = 62
"000111110",  -- sqrt(3795) = 62
"000111110",  -- sqrt(3796) = 62
"000111110",  -- sqrt(3797) = 62
"000111110",  -- sqrt(3798) = 62
"000111110",  -- sqrt(3799) = 62
"000111110",  -- sqrt(3800) = 62
"000111110",  -- sqrt(3801) = 62
"000111110",  -- sqrt(3802) = 62
"000111110",  -- sqrt(3803) = 62
"000111110",  -- sqrt(3804) = 62
"000111110",  -- sqrt(3805) = 62
"000111110",  -- sqrt(3806) = 62
"000111110",  -- sqrt(3807) = 62
"000111110",  -- sqrt(3808) = 62
"000111110",  -- sqrt(3809) = 62
"000111110",  -- sqrt(3810) = 62
"000111110",  -- sqrt(3811) = 62
"000111110",  -- sqrt(3812) = 62
"000111110",  -- sqrt(3813) = 62
"000111110",  -- sqrt(3814) = 62
"000111110",  -- sqrt(3815) = 62
"000111110",  -- sqrt(3816) = 62
"000111110",  -- sqrt(3817) = 62
"000111110",  -- sqrt(3818) = 62
"000111110",  -- sqrt(3819) = 62
"000111110",  -- sqrt(3820) = 62
"000111110",  -- sqrt(3821) = 62
"000111110",  -- sqrt(3822) = 62
"000111110",  -- sqrt(3823) = 62
"000111110",  -- sqrt(3824) = 62
"000111110",  -- sqrt(3825) = 62
"000111110",  -- sqrt(3826) = 62
"000111110",  -- sqrt(3827) = 62
"000111110",  -- sqrt(3828) = 62
"000111110",  -- sqrt(3829) = 62
"000111110",  -- sqrt(3830) = 62
"000111110",  -- sqrt(3831) = 62
"000111110",  -- sqrt(3832) = 62
"000111110",  -- sqrt(3833) = 62
"000111110",  -- sqrt(3834) = 62
"000111110",  -- sqrt(3835) = 62
"000111110",  -- sqrt(3836) = 62
"000111110",  -- sqrt(3837) = 62
"000111110",  -- sqrt(3838) = 62
"000111110",  -- sqrt(3839) = 62
"000111110",  -- sqrt(3840) = 62
"000111110",  -- sqrt(3841) = 62
"000111110",  -- sqrt(3842) = 62
"000111110",  -- sqrt(3843) = 62
"000111110",  -- sqrt(3844) = 62
"000111110",  -- sqrt(3845) = 62
"000111110",  -- sqrt(3846) = 62
"000111110",  -- sqrt(3847) = 62
"000111110",  -- sqrt(3848) = 62
"000111110",  -- sqrt(3849) = 62
"000111110",  -- sqrt(3850) = 62
"000111110",  -- sqrt(3851) = 62
"000111110",  -- sqrt(3852) = 62
"000111110",  -- sqrt(3853) = 62
"000111110",  -- sqrt(3854) = 62
"000111110",  -- sqrt(3855) = 62
"000111110",  -- sqrt(3856) = 62
"000111110",  -- sqrt(3857) = 62
"000111110",  -- sqrt(3858) = 62
"000111110",  -- sqrt(3859) = 62
"000111110",  -- sqrt(3860) = 62
"000111110",  -- sqrt(3861) = 62
"000111110",  -- sqrt(3862) = 62
"000111110",  -- sqrt(3863) = 62
"000111110",  -- sqrt(3864) = 62
"000111110",  -- sqrt(3865) = 62
"000111110",  -- sqrt(3866) = 62
"000111110",  -- sqrt(3867) = 62
"000111110",  -- sqrt(3868) = 62
"000111110",  -- sqrt(3869) = 62
"000111110",  -- sqrt(3870) = 62
"000111110",  -- sqrt(3871) = 62
"000111110",  -- sqrt(3872) = 62
"000111110",  -- sqrt(3873) = 62
"000111110",  -- sqrt(3874) = 62
"000111110",  -- sqrt(3875) = 62
"000111110",  -- sqrt(3876) = 62
"000111110",  -- sqrt(3877) = 62
"000111110",  -- sqrt(3878) = 62
"000111110",  -- sqrt(3879) = 62
"000111110",  -- sqrt(3880) = 62
"000111110",  -- sqrt(3881) = 62
"000111110",  -- sqrt(3882) = 62
"000111110",  -- sqrt(3883) = 62
"000111110",  -- sqrt(3884) = 62
"000111110",  -- sqrt(3885) = 62
"000111110",  -- sqrt(3886) = 62
"000111110",  -- sqrt(3887) = 62
"000111110",  -- sqrt(3888) = 62
"000111110",  -- sqrt(3889) = 62
"000111110",  -- sqrt(3890) = 62
"000111110",  -- sqrt(3891) = 62
"000111110",  -- sqrt(3892) = 62
"000111110",  -- sqrt(3893) = 62
"000111110",  -- sqrt(3894) = 62
"000111110",  -- sqrt(3895) = 62
"000111110",  -- sqrt(3896) = 62
"000111110",  -- sqrt(3897) = 62
"000111110",  -- sqrt(3898) = 62
"000111110",  -- sqrt(3899) = 62
"000111110",  -- sqrt(3900) = 62
"000111110",  -- sqrt(3901) = 62
"000111110",  -- sqrt(3902) = 62
"000111110",  -- sqrt(3903) = 62
"000111110",  -- sqrt(3904) = 62
"000111110",  -- sqrt(3905) = 62
"000111110",  -- sqrt(3906) = 62
"000111111",  -- sqrt(3907) = 63
"000111111",  -- sqrt(3908) = 63
"000111111",  -- sqrt(3909) = 63
"000111111",  -- sqrt(3910) = 63
"000111111",  -- sqrt(3911) = 63
"000111111",  -- sqrt(3912) = 63
"000111111",  -- sqrt(3913) = 63
"000111111",  -- sqrt(3914) = 63
"000111111",  -- sqrt(3915) = 63
"000111111",  -- sqrt(3916) = 63
"000111111",  -- sqrt(3917) = 63
"000111111",  -- sqrt(3918) = 63
"000111111",  -- sqrt(3919) = 63
"000111111",  -- sqrt(3920) = 63
"000111111",  -- sqrt(3921) = 63
"000111111",  -- sqrt(3922) = 63
"000111111",  -- sqrt(3923) = 63
"000111111",  -- sqrt(3924) = 63
"000111111",  -- sqrt(3925) = 63
"000111111",  -- sqrt(3926) = 63
"000111111",  -- sqrt(3927) = 63
"000111111",  -- sqrt(3928) = 63
"000111111",  -- sqrt(3929) = 63
"000111111",  -- sqrt(3930) = 63
"000111111",  -- sqrt(3931) = 63
"000111111",  -- sqrt(3932) = 63
"000111111",  -- sqrt(3933) = 63
"000111111",  -- sqrt(3934) = 63
"000111111",  -- sqrt(3935) = 63
"000111111",  -- sqrt(3936) = 63
"000111111",  -- sqrt(3937) = 63
"000111111",  -- sqrt(3938) = 63
"000111111",  -- sqrt(3939) = 63
"000111111",  -- sqrt(3940) = 63
"000111111",  -- sqrt(3941) = 63
"000111111",  -- sqrt(3942) = 63
"000111111",  -- sqrt(3943) = 63
"000111111",  -- sqrt(3944) = 63
"000111111",  -- sqrt(3945) = 63
"000111111",  -- sqrt(3946) = 63
"000111111",  -- sqrt(3947) = 63
"000111111",  -- sqrt(3948) = 63
"000111111",  -- sqrt(3949) = 63
"000111111",  -- sqrt(3950) = 63
"000111111",  -- sqrt(3951) = 63
"000111111",  -- sqrt(3952) = 63
"000111111",  -- sqrt(3953) = 63
"000111111",  -- sqrt(3954) = 63
"000111111",  -- sqrt(3955) = 63
"000111111",  -- sqrt(3956) = 63
"000111111",  -- sqrt(3957) = 63
"000111111",  -- sqrt(3958) = 63
"000111111",  -- sqrt(3959) = 63
"000111111",  -- sqrt(3960) = 63
"000111111",  -- sqrt(3961) = 63
"000111111",  -- sqrt(3962) = 63
"000111111",  -- sqrt(3963) = 63
"000111111",  -- sqrt(3964) = 63
"000111111",  -- sqrt(3965) = 63
"000111111",  -- sqrt(3966) = 63
"000111111",  -- sqrt(3967) = 63
"000111111",  -- sqrt(3968) = 63
"000111111",  -- sqrt(3969) = 63
"000111111",  -- sqrt(3970) = 63
"000111111",  -- sqrt(3971) = 63
"000111111",  -- sqrt(3972) = 63
"000111111",  -- sqrt(3973) = 63
"000111111",  -- sqrt(3974) = 63
"000111111",  -- sqrt(3975) = 63
"000111111",  -- sqrt(3976) = 63
"000111111",  -- sqrt(3977) = 63
"000111111",  -- sqrt(3978) = 63
"000111111",  -- sqrt(3979) = 63
"000111111",  -- sqrt(3980) = 63
"000111111",  -- sqrt(3981) = 63
"000111111",  -- sqrt(3982) = 63
"000111111",  -- sqrt(3983) = 63
"000111111",  -- sqrt(3984) = 63
"000111111",  -- sqrt(3985) = 63
"000111111",  -- sqrt(3986) = 63
"000111111",  -- sqrt(3987) = 63
"000111111",  -- sqrt(3988) = 63
"000111111",  -- sqrt(3989) = 63
"000111111",  -- sqrt(3990) = 63
"000111111",  -- sqrt(3991) = 63
"000111111",  -- sqrt(3992) = 63
"000111111",  -- sqrt(3993) = 63
"000111111",  -- sqrt(3994) = 63
"000111111",  -- sqrt(3995) = 63
"000111111",  -- sqrt(3996) = 63
"000111111",  -- sqrt(3997) = 63
"000111111",  -- sqrt(3998) = 63
"000111111",  -- sqrt(3999) = 63
"000111111",  -- sqrt(4000) = 63
"000111111",  -- sqrt(4001) = 63
"000111111",  -- sqrt(4002) = 63
"000111111",  -- sqrt(4003) = 63
"000111111",  -- sqrt(4004) = 63
"000111111",  -- sqrt(4005) = 63
"000111111",  -- sqrt(4006) = 63
"000111111",  -- sqrt(4007) = 63
"000111111",  -- sqrt(4008) = 63
"000111111",  -- sqrt(4009) = 63
"000111111",  -- sqrt(4010) = 63
"000111111",  -- sqrt(4011) = 63
"000111111",  -- sqrt(4012) = 63
"000111111",  -- sqrt(4013) = 63
"000111111",  -- sqrt(4014) = 63
"000111111",  -- sqrt(4015) = 63
"000111111",  -- sqrt(4016) = 63
"000111111",  -- sqrt(4017) = 63
"000111111",  -- sqrt(4018) = 63
"000111111",  -- sqrt(4019) = 63
"000111111",  -- sqrt(4020) = 63
"000111111",  -- sqrt(4021) = 63
"000111111",  -- sqrt(4022) = 63
"000111111",  -- sqrt(4023) = 63
"000111111",  -- sqrt(4024) = 63
"000111111",  -- sqrt(4025) = 63
"000111111",  -- sqrt(4026) = 63
"000111111",  -- sqrt(4027) = 63
"000111111",  -- sqrt(4028) = 63
"000111111",  -- sqrt(4029) = 63
"000111111",  -- sqrt(4030) = 63
"000111111",  -- sqrt(4031) = 63
"000111111",  -- sqrt(4032) = 63
"001000000",  -- sqrt(4033) = 64
"001000000",  -- sqrt(4034) = 64
"001000000",  -- sqrt(4035) = 64
"001000000",  -- sqrt(4036) = 64
"001000000",  -- sqrt(4037) = 64
"001000000",  -- sqrt(4038) = 64
"001000000",  -- sqrt(4039) = 64
"001000000",  -- sqrt(4040) = 64
"001000000",  -- sqrt(4041) = 64
"001000000",  -- sqrt(4042) = 64
"001000000",  -- sqrt(4043) = 64
"001000000",  -- sqrt(4044) = 64
"001000000",  -- sqrt(4045) = 64
"001000000",  -- sqrt(4046) = 64
"001000000",  -- sqrt(4047) = 64
"001000000",  -- sqrt(4048) = 64
"001000000",  -- sqrt(4049) = 64
"001000000",  -- sqrt(4050) = 64
"001000000",  -- sqrt(4051) = 64
"001000000",  -- sqrt(4052) = 64
"001000000",  -- sqrt(4053) = 64
"001000000",  -- sqrt(4054) = 64
"001000000",  -- sqrt(4055) = 64
"001000000",  -- sqrt(4056) = 64
"001000000",  -- sqrt(4057) = 64
"001000000",  -- sqrt(4058) = 64
"001000000",  -- sqrt(4059) = 64
"001000000",  -- sqrt(4060) = 64
"001000000",  -- sqrt(4061) = 64
"001000000",  -- sqrt(4062) = 64
"001000000",  -- sqrt(4063) = 64
"001000000",  -- sqrt(4064) = 64
"001000000",  -- sqrt(4065) = 64
"001000000",  -- sqrt(4066) = 64
"001000000",  -- sqrt(4067) = 64
"001000000",  -- sqrt(4068) = 64
"001000000",  -- sqrt(4069) = 64
"001000000",  -- sqrt(4070) = 64
"001000000",  -- sqrt(4071) = 64
"001000000",  -- sqrt(4072) = 64
"001000000",  -- sqrt(4073) = 64
"001000000",  -- sqrt(4074) = 64
"001000000",  -- sqrt(4075) = 64
"001000000",  -- sqrt(4076) = 64
"001000000",  -- sqrt(4077) = 64
"001000000",  -- sqrt(4078) = 64
"001000000",  -- sqrt(4079) = 64
"001000000",  -- sqrt(4080) = 64
"001000000",  -- sqrt(4081) = 64
"001000000",  -- sqrt(4082) = 64
"001000000",  -- sqrt(4083) = 64
"001000000",  -- sqrt(4084) = 64
"001000000",  -- sqrt(4085) = 64
"001000000",  -- sqrt(4086) = 64
"001000000",  -- sqrt(4087) = 64
"001000000",  -- sqrt(4088) = 64
"001000000",  -- sqrt(4089) = 64
"001000000",  -- sqrt(4090) = 64
"001000000",  -- sqrt(4091) = 64
"001000000",  -- sqrt(4092) = 64
"001000000",  -- sqrt(4093) = 64
"001000000",  -- sqrt(4094) = 64
"001000000",  -- sqrt(4095) = 64
"001000000",  -- sqrt(4096) = 64
"001000000",  -- sqrt(4097) = 64
"001000000",  -- sqrt(4098) = 64
"001000000",  -- sqrt(4099) = 64
"001000000",  -- sqrt(4100) = 64
"001000000",  -- sqrt(4101) = 64
"001000000",  -- sqrt(4102) = 64
"001000000",  -- sqrt(4103) = 64
"001000000",  -- sqrt(4104) = 64
"001000000",  -- sqrt(4105) = 64
"001000000",  -- sqrt(4106) = 64
"001000000",  -- sqrt(4107) = 64
"001000000",  -- sqrt(4108) = 64
"001000000",  -- sqrt(4109) = 64
"001000000",  -- sqrt(4110) = 64
"001000000",  -- sqrt(4111) = 64
"001000000",  -- sqrt(4112) = 64
"001000000",  -- sqrt(4113) = 64
"001000000",  -- sqrt(4114) = 64
"001000000",  -- sqrt(4115) = 64
"001000000",  -- sqrt(4116) = 64
"001000000",  -- sqrt(4117) = 64
"001000000",  -- sqrt(4118) = 64
"001000000",  -- sqrt(4119) = 64
"001000000",  -- sqrt(4120) = 64
"001000000",  -- sqrt(4121) = 64
"001000000",  -- sqrt(4122) = 64
"001000000",  -- sqrt(4123) = 64
"001000000",  -- sqrt(4124) = 64
"001000000",  -- sqrt(4125) = 64
"001000000",  -- sqrt(4126) = 64
"001000000",  -- sqrt(4127) = 64
"001000000",  -- sqrt(4128) = 64
"001000000",  -- sqrt(4129) = 64
"001000000",  -- sqrt(4130) = 64
"001000000",  -- sqrt(4131) = 64
"001000000",  -- sqrt(4132) = 64
"001000000",  -- sqrt(4133) = 64
"001000000",  -- sqrt(4134) = 64
"001000000",  -- sqrt(4135) = 64
"001000000",  -- sqrt(4136) = 64
"001000000",  -- sqrt(4137) = 64
"001000000",  -- sqrt(4138) = 64
"001000000",  -- sqrt(4139) = 64
"001000000",  -- sqrt(4140) = 64
"001000000",  -- sqrt(4141) = 64
"001000000",  -- sqrt(4142) = 64
"001000000",  -- sqrt(4143) = 64
"001000000",  -- sqrt(4144) = 64
"001000000",  -- sqrt(4145) = 64
"001000000",  -- sqrt(4146) = 64
"001000000",  -- sqrt(4147) = 64
"001000000",  -- sqrt(4148) = 64
"001000000",  -- sqrt(4149) = 64
"001000000",  -- sqrt(4150) = 64
"001000000",  -- sqrt(4151) = 64
"001000000",  -- sqrt(4152) = 64
"001000000",  -- sqrt(4153) = 64
"001000000",  -- sqrt(4154) = 64
"001000000",  -- sqrt(4155) = 64
"001000000",  -- sqrt(4156) = 64
"001000000",  -- sqrt(4157) = 64
"001000000",  -- sqrt(4158) = 64
"001000000",  -- sqrt(4159) = 64
"001000000",  -- sqrt(4160) = 64
"001000001",  -- sqrt(4161) = 65
"001000001",  -- sqrt(4162) = 65
"001000001",  -- sqrt(4163) = 65
"001000001",  -- sqrt(4164) = 65
"001000001",  -- sqrt(4165) = 65
"001000001",  -- sqrt(4166) = 65
"001000001",  -- sqrt(4167) = 65
"001000001",  -- sqrt(4168) = 65
"001000001",  -- sqrt(4169) = 65
"001000001",  -- sqrt(4170) = 65
"001000001",  -- sqrt(4171) = 65
"001000001",  -- sqrt(4172) = 65
"001000001",  -- sqrt(4173) = 65
"001000001",  -- sqrt(4174) = 65
"001000001",  -- sqrt(4175) = 65
"001000001",  -- sqrt(4176) = 65
"001000001",  -- sqrt(4177) = 65
"001000001",  -- sqrt(4178) = 65
"001000001",  -- sqrt(4179) = 65
"001000001",  -- sqrt(4180) = 65
"001000001",  -- sqrt(4181) = 65
"001000001",  -- sqrt(4182) = 65
"001000001",  -- sqrt(4183) = 65
"001000001",  -- sqrt(4184) = 65
"001000001",  -- sqrt(4185) = 65
"001000001",  -- sqrt(4186) = 65
"001000001",  -- sqrt(4187) = 65
"001000001",  -- sqrt(4188) = 65
"001000001",  -- sqrt(4189) = 65
"001000001",  -- sqrt(4190) = 65
"001000001",  -- sqrt(4191) = 65
"001000001",  -- sqrt(4192) = 65
"001000001",  -- sqrt(4193) = 65
"001000001",  -- sqrt(4194) = 65
"001000001",  -- sqrt(4195) = 65
"001000001",  -- sqrt(4196) = 65
"001000001",  -- sqrt(4197) = 65
"001000001",  -- sqrt(4198) = 65
"001000001",  -- sqrt(4199) = 65
"001000001",  -- sqrt(4200) = 65
"001000001",  -- sqrt(4201) = 65
"001000001",  -- sqrt(4202) = 65
"001000001",  -- sqrt(4203) = 65
"001000001",  -- sqrt(4204) = 65
"001000001",  -- sqrt(4205) = 65
"001000001",  -- sqrt(4206) = 65
"001000001",  -- sqrt(4207) = 65
"001000001",  -- sqrt(4208) = 65
"001000001",  -- sqrt(4209) = 65
"001000001",  -- sqrt(4210) = 65
"001000001",  -- sqrt(4211) = 65
"001000001",  -- sqrt(4212) = 65
"001000001",  -- sqrt(4213) = 65
"001000001",  -- sqrt(4214) = 65
"001000001",  -- sqrt(4215) = 65
"001000001",  -- sqrt(4216) = 65
"001000001",  -- sqrt(4217) = 65
"001000001",  -- sqrt(4218) = 65
"001000001",  -- sqrt(4219) = 65
"001000001",  -- sqrt(4220) = 65
"001000001",  -- sqrt(4221) = 65
"001000001",  -- sqrt(4222) = 65
"001000001",  -- sqrt(4223) = 65
"001000001",  -- sqrt(4224) = 65
"001000001",  -- sqrt(4225) = 65
"001000001",  -- sqrt(4226) = 65
"001000001",  -- sqrt(4227) = 65
"001000001",  -- sqrt(4228) = 65
"001000001",  -- sqrt(4229) = 65
"001000001",  -- sqrt(4230) = 65
"001000001",  -- sqrt(4231) = 65
"001000001",  -- sqrt(4232) = 65
"001000001",  -- sqrt(4233) = 65
"001000001",  -- sqrt(4234) = 65
"001000001",  -- sqrt(4235) = 65
"001000001",  -- sqrt(4236) = 65
"001000001",  -- sqrt(4237) = 65
"001000001",  -- sqrt(4238) = 65
"001000001",  -- sqrt(4239) = 65
"001000001",  -- sqrt(4240) = 65
"001000001",  -- sqrt(4241) = 65
"001000001",  -- sqrt(4242) = 65
"001000001",  -- sqrt(4243) = 65
"001000001",  -- sqrt(4244) = 65
"001000001",  -- sqrt(4245) = 65
"001000001",  -- sqrt(4246) = 65
"001000001",  -- sqrt(4247) = 65
"001000001",  -- sqrt(4248) = 65
"001000001",  -- sqrt(4249) = 65
"001000001",  -- sqrt(4250) = 65
"001000001",  -- sqrt(4251) = 65
"001000001",  -- sqrt(4252) = 65
"001000001",  -- sqrt(4253) = 65
"001000001",  -- sqrt(4254) = 65
"001000001",  -- sqrt(4255) = 65
"001000001",  -- sqrt(4256) = 65
"001000001",  -- sqrt(4257) = 65
"001000001",  -- sqrt(4258) = 65
"001000001",  -- sqrt(4259) = 65
"001000001",  -- sqrt(4260) = 65
"001000001",  -- sqrt(4261) = 65
"001000001",  -- sqrt(4262) = 65
"001000001",  -- sqrt(4263) = 65
"001000001",  -- sqrt(4264) = 65
"001000001",  -- sqrt(4265) = 65
"001000001",  -- sqrt(4266) = 65
"001000001",  -- sqrt(4267) = 65
"001000001",  -- sqrt(4268) = 65
"001000001",  -- sqrt(4269) = 65
"001000001",  -- sqrt(4270) = 65
"001000001",  -- sqrt(4271) = 65
"001000001",  -- sqrt(4272) = 65
"001000001",  -- sqrt(4273) = 65
"001000001",  -- sqrt(4274) = 65
"001000001",  -- sqrt(4275) = 65
"001000001",  -- sqrt(4276) = 65
"001000001",  -- sqrt(4277) = 65
"001000001",  -- sqrt(4278) = 65
"001000001",  -- sqrt(4279) = 65
"001000001",  -- sqrt(4280) = 65
"001000001",  -- sqrt(4281) = 65
"001000001",  -- sqrt(4282) = 65
"001000001",  -- sqrt(4283) = 65
"001000001",  -- sqrt(4284) = 65
"001000001",  -- sqrt(4285) = 65
"001000001",  -- sqrt(4286) = 65
"001000001",  -- sqrt(4287) = 65
"001000001",  -- sqrt(4288) = 65
"001000001",  -- sqrt(4289) = 65
"001000001",  -- sqrt(4290) = 65
"001000010",  -- sqrt(4291) = 66
"001000010",  -- sqrt(4292) = 66
"001000010",  -- sqrt(4293) = 66
"001000010",  -- sqrt(4294) = 66
"001000010",  -- sqrt(4295) = 66
"001000010",  -- sqrt(4296) = 66
"001000010",  -- sqrt(4297) = 66
"001000010",  -- sqrt(4298) = 66
"001000010",  -- sqrt(4299) = 66
"001000010",  -- sqrt(4300) = 66
"001000010",  -- sqrt(4301) = 66
"001000010",  -- sqrt(4302) = 66
"001000010",  -- sqrt(4303) = 66
"001000010",  -- sqrt(4304) = 66
"001000010",  -- sqrt(4305) = 66
"001000010",  -- sqrt(4306) = 66
"001000010",  -- sqrt(4307) = 66
"001000010",  -- sqrt(4308) = 66
"001000010",  -- sqrt(4309) = 66
"001000010",  -- sqrt(4310) = 66
"001000010",  -- sqrt(4311) = 66
"001000010",  -- sqrt(4312) = 66
"001000010",  -- sqrt(4313) = 66
"001000010",  -- sqrt(4314) = 66
"001000010",  -- sqrt(4315) = 66
"001000010",  -- sqrt(4316) = 66
"001000010",  -- sqrt(4317) = 66
"001000010",  -- sqrt(4318) = 66
"001000010",  -- sqrt(4319) = 66
"001000010",  -- sqrt(4320) = 66
"001000010",  -- sqrt(4321) = 66
"001000010",  -- sqrt(4322) = 66
"001000010",  -- sqrt(4323) = 66
"001000010",  -- sqrt(4324) = 66
"001000010",  -- sqrt(4325) = 66
"001000010",  -- sqrt(4326) = 66
"001000010",  -- sqrt(4327) = 66
"001000010",  -- sqrt(4328) = 66
"001000010",  -- sqrt(4329) = 66
"001000010",  -- sqrt(4330) = 66
"001000010",  -- sqrt(4331) = 66
"001000010",  -- sqrt(4332) = 66
"001000010",  -- sqrt(4333) = 66
"001000010",  -- sqrt(4334) = 66
"001000010",  -- sqrt(4335) = 66
"001000010",  -- sqrt(4336) = 66
"001000010",  -- sqrt(4337) = 66
"001000010",  -- sqrt(4338) = 66
"001000010",  -- sqrt(4339) = 66
"001000010",  -- sqrt(4340) = 66
"001000010",  -- sqrt(4341) = 66
"001000010",  -- sqrt(4342) = 66
"001000010",  -- sqrt(4343) = 66
"001000010",  -- sqrt(4344) = 66
"001000010",  -- sqrt(4345) = 66
"001000010",  -- sqrt(4346) = 66
"001000010",  -- sqrt(4347) = 66
"001000010",  -- sqrt(4348) = 66
"001000010",  -- sqrt(4349) = 66
"001000010",  -- sqrt(4350) = 66
"001000010",  -- sqrt(4351) = 66
"001000010",  -- sqrt(4352) = 66
"001000010",  -- sqrt(4353) = 66
"001000010",  -- sqrt(4354) = 66
"001000010",  -- sqrt(4355) = 66
"001000010",  -- sqrt(4356) = 66
"001000010",  -- sqrt(4357) = 66
"001000010",  -- sqrt(4358) = 66
"001000010",  -- sqrt(4359) = 66
"001000010",  -- sqrt(4360) = 66
"001000010",  -- sqrt(4361) = 66
"001000010",  -- sqrt(4362) = 66
"001000010",  -- sqrt(4363) = 66
"001000010",  -- sqrt(4364) = 66
"001000010",  -- sqrt(4365) = 66
"001000010",  -- sqrt(4366) = 66
"001000010",  -- sqrt(4367) = 66
"001000010",  -- sqrt(4368) = 66
"001000010",  -- sqrt(4369) = 66
"001000010",  -- sqrt(4370) = 66
"001000010",  -- sqrt(4371) = 66
"001000010",  -- sqrt(4372) = 66
"001000010",  -- sqrt(4373) = 66
"001000010",  -- sqrt(4374) = 66
"001000010",  -- sqrt(4375) = 66
"001000010",  -- sqrt(4376) = 66
"001000010",  -- sqrt(4377) = 66
"001000010",  -- sqrt(4378) = 66
"001000010",  -- sqrt(4379) = 66
"001000010",  -- sqrt(4380) = 66
"001000010",  -- sqrt(4381) = 66
"001000010",  -- sqrt(4382) = 66
"001000010",  -- sqrt(4383) = 66
"001000010",  -- sqrt(4384) = 66
"001000010",  -- sqrt(4385) = 66
"001000010",  -- sqrt(4386) = 66
"001000010",  -- sqrt(4387) = 66
"001000010",  -- sqrt(4388) = 66
"001000010",  -- sqrt(4389) = 66
"001000010",  -- sqrt(4390) = 66
"001000010",  -- sqrt(4391) = 66
"001000010",  -- sqrt(4392) = 66
"001000010",  -- sqrt(4393) = 66
"001000010",  -- sqrt(4394) = 66
"001000010",  -- sqrt(4395) = 66
"001000010",  -- sqrt(4396) = 66
"001000010",  -- sqrt(4397) = 66
"001000010",  -- sqrt(4398) = 66
"001000010",  -- sqrt(4399) = 66
"001000010",  -- sqrt(4400) = 66
"001000010",  -- sqrt(4401) = 66
"001000010",  -- sqrt(4402) = 66
"001000010",  -- sqrt(4403) = 66
"001000010",  -- sqrt(4404) = 66
"001000010",  -- sqrt(4405) = 66
"001000010",  -- sqrt(4406) = 66
"001000010",  -- sqrt(4407) = 66
"001000010",  -- sqrt(4408) = 66
"001000010",  -- sqrt(4409) = 66
"001000010",  -- sqrt(4410) = 66
"001000010",  -- sqrt(4411) = 66
"001000010",  -- sqrt(4412) = 66
"001000010",  -- sqrt(4413) = 66
"001000010",  -- sqrt(4414) = 66
"001000010",  -- sqrt(4415) = 66
"001000010",  -- sqrt(4416) = 66
"001000010",  -- sqrt(4417) = 66
"001000010",  -- sqrt(4418) = 66
"001000010",  -- sqrt(4419) = 66
"001000010",  -- sqrt(4420) = 66
"001000010",  -- sqrt(4421) = 66
"001000010",  -- sqrt(4422) = 66
"001000011",  -- sqrt(4423) = 67
"001000011",  -- sqrt(4424) = 67
"001000011",  -- sqrt(4425) = 67
"001000011",  -- sqrt(4426) = 67
"001000011",  -- sqrt(4427) = 67
"001000011",  -- sqrt(4428) = 67
"001000011",  -- sqrt(4429) = 67
"001000011",  -- sqrt(4430) = 67
"001000011",  -- sqrt(4431) = 67
"001000011",  -- sqrt(4432) = 67
"001000011",  -- sqrt(4433) = 67
"001000011",  -- sqrt(4434) = 67
"001000011",  -- sqrt(4435) = 67
"001000011",  -- sqrt(4436) = 67
"001000011",  -- sqrt(4437) = 67
"001000011",  -- sqrt(4438) = 67
"001000011",  -- sqrt(4439) = 67
"001000011",  -- sqrt(4440) = 67
"001000011",  -- sqrt(4441) = 67
"001000011",  -- sqrt(4442) = 67
"001000011",  -- sqrt(4443) = 67
"001000011",  -- sqrt(4444) = 67
"001000011",  -- sqrt(4445) = 67
"001000011",  -- sqrt(4446) = 67
"001000011",  -- sqrt(4447) = 67
"001000011",  -- sqrt(4448) = 67
"001000011",  -- sqrt(4449) = 67
"001000011",  -- sqrt(4450) = 67
"001000011",  -- sqrt(4451) = 67
"001000011",  -- sqrt(4452) = 67
"001000011",  -- sqrt(4453) = 67
"001000011",  -- sqrt(4454) = 67
"001000011",  -- sqrt(4455) = 67
"001000011",  -- sqrt(4456) = 67
"001000011",  -- sqrt(4457) = 67
"001000011",  -- sqrt(4458) = 67
"001000011",  -- sqrt(4459) = 67
"001000011",  -- sqrt(4460) = 67
"001000011",  -- sqrt(4461) = 67
"001000011",  -- sqrt(4462) = 67
"001000011",  -- sqrt(4463) = 67
"001000011",  -- sqrt(4464) = 67
"001000011",  -- sqrt(4465) = 67
"001000011",  -- sqrt(4466) = 67
"001000011",  -- sqrt(4467) = 67
"001000011",  -- sqrt(4468) = 67
"001000011",  -- sqrt(4469) = 67
"001000011",  -- sqrt(4470) = 67
"001000011",  -- sqrt(4471) = 67
"001000011",  -- sqrt(4472) = 67
"001000011",  -- sqrt(4473) = 67
"001000011",  -- sqrt(4474) = 67
"001000011",  -- sqrt(4475) = 67
"001000011",  -- sqrt(4476) = 67
"001000011",  -- sqrt(4477) = 67
"001000011",  -- sqrt(4478) = 67
"001000011",  -- sqrt(4479) = 67
"001000011",  -- sqrt(4480) = 67
"001000011",  -- sqrt(4481) = 67
"001000011",  -- sqrt(4482) = 67
"001000011",  -- sqrt(4483) = 67
"001000011",  -- sqrt(4484) = 67
"001000011",  -- sqrt(4485) = 67
"001000011",  -- sqrt(4486) = 67
"001000011",  -- sqrt(4487) = 67
"001000011",  -- sqrt(4488) = 67
"001000011",  -- sqrt(4489) = 67
"001000011",  -- sqrt(4490) = 67
"001000011",  -- sqrt(4491) = 67
"001000011",  -- sqrt(4492) = 67
"001000011",  -- sqrt(4493) = 67
"001000011",  -- sqrt(4494) = 67
"001000011",  -- sqrt(4495) = 67
"001000011",  -- sqrt(4496) = 67
"001000011",  -- sqrt(4497) = 67
"001000011",  -- sqrt(4498) = 67
"001000011",  -- sqrt(4499) = 67
"001000011",  -- sqrt(4500) = 67
"001000011",  -- sqrt(4501) = 67
"001000011",  -- sqrt(4502) = 67
"001000011",  -- sqrt(4503) = 67
"001000011",  -- sqrt(4504) = 67
"001000011",  -- sqrt(4505) = 67
"001000011",  -- sqrt(4506) = 67
"001000011",  -- sqrt(4507) = 67
"001000011",  -- sqrt(4508) = 67
"001000011",  -- sqrt(4509) = 67
"001000011",  -- sqrt(4510) = 67
"001000011",  -- sqrt(4511) = 67
"001000011",  -- sqrt(4512) = 67
"001000011",  -- sqrt(4513) = 67
"001000011",  -- sqrt(4514) = 67
"001000011",  -- sqrt(4515) = 67
"001000011",  -- sqrt(4516) = 67
"001000011",  -- sqrt(4517) = 67
"001000011",  -- sqrt(4518) = 67
"001000011",  -- sqrt(4519) = 67
"001000011",  -- sqrt(4520) = 67
"001000011",  -- sqrt(4521) = 67
"001000011",  -- sqrt(4522) = 67
"001000011",  -- sqrt(4523) = 67
"001000011",  -- sqrt(4524) = 67
"001000011",  -- sqrt(4525) = 67
"001000011",  -- sqrt(4526) = 67
"001000011",  -- sqrt(4527) = 67
"001000011",  -- sqrt(4528) = 67
"001000011",  -- sqrt(4529) = 67
"001000011",  -- sqrt(4530) = 67
"001000011",  -- sqrt(4531) = 67
"001000011",  -- sqrt(4532) = 67
"001000011",  -- sqrt(4533) = 67
"001000011",  -- sqrt(4534) = 67
"001000011",  -- sqrt(4535) = 67
"001000011",  -- sqrt(4536) = 67
"001000011",  -- sqrt(4537) = 67
"001000011",  -- sqrt(4538) = 67
"001000011",  -- sqrt(4539) = 67
"001000011",  -- sqrt(4540) = 67
"001000011",  -- sqrt(4541) = 67
"001000011",  -- sqrt(4542) = 67
"001000011",  -- sqrt(4543) = 67
"001000011",  -- sqrt(4544) = 67
"001000011",  -- sqrt(4545) = 67
"001000011",  -- sqrt(4546) = 67
"001000011",  -- sqrt(4547) = 67
"001000011",  -- sqrt(4548) = 67
"001000011",  -- sqrt(4549) = 67
"001000011",  -- sqrt(4550) = 67
"001000011",  -- sqrt(4551) = 67
"001000011",  -- sqrt(4552) = 67
"001000011",  -- sqrt(4553) = 67
"001000011",  -- sqrt(4554) = 67
"001000011",  -- sqrt(4555) = 67
"001000011",  -- sqrt(4556) = 67
"001000100",  -- sqrt(4557) = 68
"001000100",  -- sqrt(4558) = 68
"001000100",  -- sqrt(4559) = 68
"001000100",  -- sqrt(4560) = 68
"001000100",  -- sqrt(4561) = 68
"001000100",  -- sqrt(4562) = 68
"001000100",  -- sqrt(4563) = 68
"001000100",  -- sqrt(4564) = 68
"001000100",  -- sqrt(4565) = 68
"001000100",  -- sqrt(4566) = 68
"001000100",  -- sqrt(4567) = 68
"001000100",  -- sqrt(4568) = 68
"001000100",  -- sqrt(4569) = 68
"001000100",  -- sqrt(4570) = 68
"001000100",  -- sqrt(4571) = 68
"001000100",  -- sqrt(4572) = 68
"001000100",  -- sqrt(4573) = 68
"001000100",  -- sqrt(4574) = 68
"001000100",  -- sqrt(4575) = 68
"001000100",  -- sqrt(4576) = 68
"001000100",  -- sqrt(4577) = 68
"001000100",  -- sqrt(4578) = 68
"001000100",  -- sqrt(4579) = 68
"001000100",  -- sqrt(4580) = 68
"001000100",  -- sqrt(4581) = 68
"001000100",  -- sqrt(4582) = 68
"001000100",  -- sqrt(4583) = 68
"001000100",  -- sqrt(4584) = 68
"001000100",  -- sqrt(4585) = 68
"001000100",  -- sqrt(4586) = 68
"001000100",  -- sqrt(4587) = 68
"001000100",  -- sqrt(4588) = 68
"001000100",  -- sqrt(4589) = 68
"001000100",  -- sqrt(4590) = 68
"001000100",  -- sqrt(4591) = 68
"001000100",  -- sqrt(4592) = 68
"001000100",  -- sqrt(4593) = 68
"001000100",  -- sqrt(4594) = 68
"001000100",  -- sqrt(4595) = 68
"001000100",  -- sqrt(4596) = 68
"001000100",  -- sqrt(4597) = 68
"001000100",  -- sqrt(4598) = 68
"001000100",  -- sqrt(4599) = 68
"001000100",  -- sqrt(4600) = 68
"001000100",  -- sqrt(4601) = 68
"001000100",  -- sqrt(4602) = 68
"001000100",  -- sqrt(4603) = 68
"001000100",  -- sqrt(4604) = 68
"001000100",  -- sqrt(4605) = 68
"001000100",  -- sqrt(4606) = 68
"001000100",  -- sqrt(4607) = 68
"001000100",  -- sqrt(4608) = 68
"001000100",  -- sqrt(4609) = 68
"001000100",  -- sqrt(4610) = 68
"001000100",  -- sqrt(4611) = 68
"001000100",  -- sqrt(4612) = 68
"001000100",  -- sqrt(4613) = 68
"001000100",  -- sqrt(4614) = 68
"001000100",  -- sqrt(4615) = 68
"001000100",  -- sqrt(4616) = 68
"001000100",  -- sqrt(4617) = 68
"001000100",  -- sqrt(4618) = 68
"001000100",  -- sqrt(4619) = 68
"001000100",  -- sqrt(4620) = 68
"001000100",  -- sqrt(4621) = 68
"001000100",  -- sqrt(4622) = 68
"001000100",  -- sqrt(4623) = 68
"001000100",  -- sqrt(4624) = 68
"001000100",  -- sqrt(4625) = 68
"001000100",  -- sqrt(4626) = 68
"001000100",  -- sqrt(4627) = 68
"001000100",  -- sqrt(4628) = 68
"001000100",  -- sqrt(4629) = 68
"001000100",  -- sqrt(4630) = 68
"001000100",  -- sqrt(4631) = 68
"001000100",  -- sqrt(4632) = 68
"001000100",  -- sqrt(4633) = 68
"001000100",  -- sqrt(4634) = 68
"001000100",  -- sqrt(4635) = 68
"001000100",  -- sqrt(4636) = 68
"001000100",  -- sqrt(4637) = 68
"001000100",  -- sqrt(4638) = 68
"001000100",  -- sqrt(4639) = 68
"001000100",  -- sqrt(4640) = 68
"001000100",  -- sqrt(4641) = 68
"001000100",  -- sqrt(4642) = 68
"001000100",  -- sqrt(4643) = 68
"001000100",  -- sqrt(4644) = 68
"001000100",  -- sqrt(4645) = 68
"001000100",  -- sqrt(4646) = 68
"001000100",  -- sqrt(4647) = 68
"001000100",  -- sqrt(4648) = 68
"001000100",  -- sqrt(4649) = 68
"001000100",  -- sqrt(4650) = 68
"001000100",  -- sqrt(4651) = 68
"001000100",  -- sqrt(4652) = 68
"001000100",  -- sqrt(4653) = 68
"001000100",  -- sqrt(4654) = 68
"001000100",  -- sqrt(4655) = 68
"001000100",  -- sqrt(4656) = 68
"001000100",  -- sqrt(4657) = 68
"001000100",  -- sqrt(4658) = 68
"001000100",  -- sqrt(4659) = 68
"001000100",  -- sqrt(4660) = 68
"001000100",  -- sqrt(4661) = 68
"001000100",  -- sqrt(4662) = 68
"001000100",  -- sqrt(4663) = 68
"001000100",  -- sqrt(4664) = 68
"001000100",  -- sqrt(4665) = 68
"001000100",  -- sqrt(4666) = 68
"001000100",  -- sqrt(4667) = 68
"001000100",  -- sqrt(4668) = 68
"001000100",  -- sqrt(4669) = 68
"001000100",  -- sqrt(4670) = 68
"001000100",  -- sqrt(4671) = 68
"001000100",  -- sqrt(4672) = 68
"001000100",  -- sqrt(4673) = 68
"001000100",  -- sqrt(4674) = 68
"001000100",  -- sqrt(4675) = 68
"001000100",  -- sqrt(4676) = 68
"001000100",  -- sqrt(4677) = 68
"001000100",  -- sqrt(4678) = 68
"001000100",  -- sqrt(4679) = 68
"001000100",  -- sqrt(4680) = 68
"001000100",  -- sqrt(4681) = 68
"001000100",  -- sqrt(4682) = 68
"001000100",  -- sqrt(4683) = 68
"001000100",  -- sqrt(4684) = 68
"001000100",  -- sqrt(4685) = 68
"001000100",  -- sqrt(4686) = 68
"001000100",  -- sqrt(4687) = 68
"001000100",  -- sqrt(4688) = 68
"001000100",  -- sqrt(4689) = 68
"001000100",  -- sqrt(4690) = 68
"001000100",  -- sqrt(4691) = 68
"001000100",  -- sqrt(4692) = 68
"001000101",  -- sqrt(4693) = 69
"001000101",  -- sqrt(4694) = 69
"001000101",  -- sqrt(4695) = 69
"001000101",  -- sqrt(4696) = 69
"001000101",  -- sqrt(4697) = 69
"001000101",  -- sqrt(4698) = 69
"001000101",  -- sqrt(4699) = 69
"001000101",  -- sqrt(4700) = 69
"001000101",  -- sqrt(4701) = 69
"001000101",  -- sqrt(4702) = 69
"001000101",  -- sqrt(4703) = 69
"001000101",  -- sqrt(4704) = 69
"001000101",  -- sqrt(4705) = 69
"001000101",  -- sqrt(4706) = 69
"001000101",  -- sqrt(4707) = 69
"001000101",  -- sqrt(4708) = 69
"001000101",  -- sqrt(4709) = 69
"001000101",  -- sqrt(4710) = 69
"001000101",  -- sqrt(4711) = 69
"001000101",  -- sqrt(4712) = 69
"001000101",  -- sqrt(4713) = 69
"001000101",  -- sqrt(4714) = 69
"001000101",  -- sqrt(4715) = 69
"001000101",  -- sqrt(4716) = 69
"001000101",  -- sqrt(4717) = 69
"001000101",  -- sqrt(4718) = 69
"001000101",  -- sqrt(4719) = 69
"001000101",  -- sqrt(4720) = 69
"001000101",  -- sqrt(4721) = 69
"001000101",  -- sqrt(4722) = 69
"001000101",  -- sqrt(4723) = 69
"001000101",  -- sqrt(4724) = 69
"001000101",  -- sqrt(4725) = 69
"001000101",  -- sqrt(4726) = 69
"001000101",  -- sqrt(4727) = 69
"001000101",  -- sqrt(4728) = 69
"001000101",  -- sqrt(4729) = 69
"001000101",  -- sqrt(4730) = 69
"001000101",  -- sqrt(4731) = 69
"001000101",  -- sqrt(4732) = 69
"001000101",  -- sqrt(4733) = 69
"001000101",  -- sqrt(4734) = 69
"001000101",  -- sqrt(4735) = 69
"001000101",  -- sqrt(4736) = 69
"001000101",  -- sqrt(4737) = 69
"001000101",  -- sqrt(4738) = 69
"001000101",  -- sqrt(4739) = 69
"001000101",  -- sqrt(4740) = 69
"001000101",  -- sqrt(4741) = 69
"001000101",  -- sqrt(4742) = 69
"001000101",  -- sqrt(4743) = 69
"001000101",  -- sqrt(4744) = 69
"001000101",  -- sqrt(4745) = 69
"001000101",  -- sqrt(4746) = 69
"001000101",  -- sqrt(4747) = 69
"001000101",  -- sqrt(4748) = 69
"001000101",  -- sqrt(4749) = 69
"001000101",  -- sqrt(4750) = 69
"001000101",  -- sqrt(4751) = 69
"001000101",  -- sqrt(4752) = 69
"001000101",  -- sqrt(4753) = 69
"001000101",  -- sqrt(4754) = 69
"001000101",  -- sqrt(4755) = 69
"001000101",  -- sqrt(4756) = 69
"001000101",  -- sqrt(4757) = 69
"001000101",  -- sqrt(4758) = 69
"001000101",  -- sqrt(4759) = 69
"001000101",  -- sqrt(4760) = 69
"001000101",  -- sqrt(4761) = 69
"001000101",  -- sqrt(4762) = 69
"001000101",  -- sqrt(4763) = 69
"001000101",  -- sqrt(4764) = 69
"001000101",  -- sqrt(4765) = 69
"001000101",  -- sqrt(4766) = 69
"001000101",  -- sqrt(4767) = 69
"001000101",  -- sqrt(4768) = 69
"001000101",  -- sqrt(4769) = 69
"001000101",  -- sqrt(4770) = 69
"001000101",  -- sqrt(4771) = 69
"001000101",  -- sqrt(4772) = 69
"001000101",  -- sqrt(4773) = 69
"001000101",  -- sqrt(4774) = 69
"001000101",  -- sqrt(4775) = 69
"001000101",  -- sqrt(4776) = 69
"001000101",  -- sqrt(4777) = 69
"001000101",  -- sqrt(4778) = 69
"001000101",  -- sqrt(4779) = 69
"001000101",  -- sqrt(4780) = 69
"001000101",  -- sqrt(4781) = 69
"001000101",  -- sqrt(4782) = 69
"001000101",  -- sqrt(4783) = 69
"001000101",  -- sqrt(4784) = 69
"001000101",  -- sqrt(4785) = 69
"001000101",  -- sqrt(4786) = 69
"001000101",  -- sqrt(4787) = 69
"001000101",  -- sqrt(4788) = 69
"001000101",  -- sqrt(4789) = 69
"001000101",  -- sqrt(4790) = 69
"001000101",  -- sqrt(4791) = 69
"001000101",  -- sqrt(4792) = 69
"001000101",  -- sqrt(4793) = 69
"001000101",  -- sqrt(4794) = 69
"001000101",  -- sqrt(4795) = 69
"001000101",  -- sqrt(4796) = 69
"001000101",  -- sqrt(4797) = 69
"001000101",  -- sqrt(4798) = 69
"001000101",  -- sqrt(4799) = 69
"001000101",  -- sqrt(4800) = 69
"001000101",  -- sqrt(4801) = 69
"001000101",  -- sqrt(4802) = 69
"001000101",  -- sqrt(4803) = 69
"001000101",  -- sqrt(4804) = 69
"001000101",  -- sqrt(4805) = 69
"001000101",  -- sqrt(4806) = 69
"001000101",  -- sqrt(4807) = 69
"001000101",  -- sqrt(4808) = 69
"001000101",  -- sqrt(4809) = 69
"001000101",  -- sqrt(4810) = 69
"001000101",  -- sqrt(4811) = 69
"001000101",  -- sqrt(4812) = 69
"001000101",  -- sqrt(4813) = 69
"001000101",  -- sqrt(4814) = 69
"001000101",  -- sqrt(4815) = 69
"001000101",  -- sqrt(4816) = 69
"001000101",  -- sqrt(4817) = 69
"001000101",  -- sqrt(4818) = 69
"001000101",  -- sqrt(4819) = 69
"001000101",  -- sqrt(4820) = 69
"001000101",  -- sqrt(4821) = 69
"001000101",  -- sqrt(4822) = 69
"001000101",  -- sqrt(4823) = 69
"001000101",  -- sqrt(4824) = 69
"001000101",  -- sqrt(4825) = 69
"001000101",  -- sqrt(4826) = 69
"001000101",  -- sqrt(4827) = 69
"001000101",  -- sqrt(4828) = 69
"001000101",  -- sqrt(4829) = 69
"001000101",  -- sqrt(4830) = 69
"001000110",  -- sqrt(4831) = 70
"001000110",  -- sqrt(4832) = 70
"001000110",  -- sqrt(4833) = 70
"001000110",  -- sqrt(4834) = 70
"001000110",  -- sqrt(4835) = 70
"001000110",  -- sqrt(4836) = 70
"001000110",  -- sqrt(4837) = 70
"001000110",  -- sqrt(4838) = 70
"001000110",  -- sqrt(4839) = 70
"001000110",  -- sqrt(4840) = 70
"001000110",  -- sqrt(4841) = 70
"001000110",  -- sqrt(4842) = 70
"001000110",  -- sqrt(4843) = 70
"001000110",  -- sqrt(4844) = 70
"001000110",  -- sqrt(4845) = 70
"001000110",  -- sqrt(4846) = 70
"001000110",  -- sqrt(4847) = 70
"001000110",  -- sqrt(4848) = 70
"001000110",  -- sqrt(4849) = 70
"001000110",  -- sqrt(4850) = 70
"001000110",  -- sqrt(4851) = 70
"001000110",  -- sqrt(4852) = 70
"001000110",  -- sqrt(4853) = 70
"001000110",  -- sqrt(4854) = 70
"001000110",  -- sqrt(4855) = 70
"001000110",  -- sqrt(4856) = 70
"001000110",  -- sqrt(4857) = 70
"001000110",  -- sqrt(4858) = 70
"001000110",  -- sqrt(4859) = 70
"001000110",  -- sqrt(4860) = 70
"001000110",  -- sqrt(4861) = 70
"001000110",  -- sqrt(4862) = 70
"001000110",  -- sqrt(4863) = 70
"001000110",  -- sqrt(4864) = 70
"001000110",  -- sqrt(4865) = 70
"001000110",  -- sqrt(4866) = 70
"001000110",  -- sqrt(4867) = 70
"001000110",  -- sqrt(4868) = 70
"001000110",  -- sqrt(4869) = 70
"001000110",  -- sqrt(4870) = 70
"001000110",  -- sqrt(4871) = 70
"001000110",  -- sqrt(4872) = 70
"001000110",  -- sqrt(4873) = 70
"001000110",  -- sqrt(4874) = 70
"001000110",  -- sqrt(4875) = 70
"001000110",  -- sqrt(4876) = 70
"001000110",  -- sqrt(4877) = 70
"001000110",  -- sqrt(4878) = 70
"001000110",  -- sqrt(4879) = 70
"001000110",  -- sqrt(4880) = 70
"001000110",  -- sqrt(4881) = 70
"001000110",  -- sqrt(4882) = 70
"001000110",  -- sqrt(4883) = 70
"001000110",  -- sqrt(4884) = 70
"001000110",  -- sqrt(4885) = 70
"001000110",  -- sqrt(4886) = 70
"001000110",  -- sqrt(4887) = 70
"001000110",  -- sqrt(4888) = 70
"001000110",  -- sqrt(4889) = 70
"001000110",  -- sqrt(4890) = 70
"001000110",  -- sqrt(4891) = 70
"001000110",  -- sqrt(4892) = 70
"001000110",  -- sqrt(4893) = 70
"001000110",  -- sqrt(4894) = 70
"001000110",  -- sqrt(4895) = 70
"001000110",  -- sqrt(4896) = 70
"001000110",  -- sqrt(4897) = 70
"001000110",  -- sqrt(4898) = 70
"001000110",  -- sqrt(4899) = 70
"001000110",  -- sqrt(4900) = 70
"001000110",  -- sqrt(4901) = 70
"001000110",  -- sqrt(4902) = 70
"001000110",  -- sqrt(4903) = 70
"001000110",  -- sqrt(4904) = 70
"001000110",  -- sqrt(4905) = 70
"001000110",  -- sqrt(4906) = 70
"001000110",  -- sqrt(4907) = 70
"001000110",  -- sqrt(4908) = 70
"001000110",  -- sqrt(4909) = 70
"001000110",  -- sqrt(4910) = 70
"001000110",  -- sqrt(4911) = 70
"001000110",  -- sqrt(4912) = 70
"001000110",  -- sqrt(4913) = 70
"001000110",  -- sqrt(4914) = 70
"001000110",  -- sqrt(4915) = 70
"001000110",  -- sqrt(4916) = 70
"001000110",  -- sqrt(4917) = 70
"001000110",  -- sqrt(4918) = 70
"001000110",  -- sqrt(4919) = 70
"001000110",  -- sqrt(4920) = 70
"001000110",  -- sqrt(4921) = 70
"001000110",  -- sqrt(4922) = 70
"001000110",  -- sqrt(4923) = 70
"001000110",  -- sqrt(4924) = 70
"001000110",  -- sqrt(4925) = 70
"001000110",  -- sqrt(4926) = 70
"001000110",  -- sqrt(4927) = 70
"001000110",  -- sqrt(4928) = 70
"001000110",  -- sqrt(4929) = 70
"001000110",  -- sqrt(4930) = 70
"001000110",  -- sqrt(4931) = 70
"001000110",  -- sqrt(4932) = 70
"001000110",  -- sqrt(4933) = 70
"001000110",  -- sqrt(4934) = 70
"001000110",  -- sqrt(4935) = 70
"001000110",  -- sqrt(4936) = 70
"001000110",  -- sqrt(4937) = 70
"001000110",  -- sqrt(4938) = 70
"001000110",  -- sqrt(4939) = 70
"001000110",  -- sqrt(4940) = 70
"001000110",  -- sqrt(4941) = 70
"001000110",  -- sqrt(4942) = 70
"001000110",  -- sqrt(4943) = 70
"001000110",  -- sqrt(4944) = 70
"001000110",  -- sqrt(4945) = 70
"001000110",  -- sqrt(4946) = 70
"001000110",  -- sqrt(4947) = 70
"001000110",  -- sqrt(4948) = 70
"001000110",  -- sqrt(4949) = 70
"001000110",  -- sqrt(4950) = 70
"001000110",  -- sqrt(4951) = 70
"001000110",  -- sqrt(4952) = 70
"001000110",  -- sqrt(4953) = 70
"001000110",  -- sqrt(4954) = 70
"001000110",  -- sqrt(4955) = 70
"001000110",  -- sqrt(4956) = 70
"001000110",  -- sqrt(4957) = 70
"001000110",  -- sqrt(4958) = 70
"001000110",  -- sqrt(4959) = 70
"001000110",  -- sqrt(4960) = 70
"001000110",  -- sqrt(4961) = 70
"001000110",  -- sqrt(4962) = 70
"001000110",  -- sqrt(4963) = 70
"001000110",  -- sqrt(4964) = 70
"001000110",  -- sqrt(4965) = 70
"001000110",  -- sqrt(4966) = 70
"001000110",  -- sqrt(4967) = 70
"001000110",  -- sqrt(4968) = 70
"001000110",  -- sqrt(4969) = 70
"001000110",  -- sqrt(4970) = 70
"001000111",  -- sqrt(4971) = 71
"001000111",  -- sqrt(4972) = 71
"001000111",  -- sqrt(4973) = 71
"001000111",  -- sqrt(4974) = 71
"001000111",  -- sqrt(4975) = 71
"001000111",  -- sqrt(4976) = 71
"001000111",  -- sqrt(4977) = 71
"001000111",  -- sqrt(4978) = 71
"001000111",  -- sqrt(4979) = 71
"001000111",  -- sqrt(4980) = 71
"001000111",  -- sqrt(4981) = 71
"001000111",  -- sqrt(4982) = 71
"001000111",  -- sqrt(4983) = 71
"001000111",  -- sqrt(4984) = 71
"001000111",  -- sqrt(4985) = 71
"001000111",  -- sqrt(4986) = 71
"001000111",  -- sqrt(4987) = 71
"001000111",  -- sqrt(4988) = 71
"001000111",  -- sqrt(4989) = 71
"001000111",  -- sqrt(4990) = 71
"001000111",  -- sqrt(4991) = 71
"001000111",  -- sqrt(4992) = 71
"001000111",  -- sqrt(4993) = 71
"001000111",  -- sqrt(4994) = 71
"001000111",  -- sqrt(4995) = 71
"001000111",  -- sqrt(4996) = 71
"001000111",  -- sqrt(4997) = 71
"001000111",  -- sqrt(4998) = 71
"001000111",  -- sqrt(4999) = 71
"001000111",  -- sqrt(5000) = 71
"001000111",  -- sqrt(5001) = 71
"001000111",  -- sqrt(5002) = 71
"001000111",  -- sqrt(5003) = 71
"001000111",  -- sqrt(5004) = 71
"001000111",  -- sqrt(5005) = 71
"001000111",  -- sqrt(5006) = 71
"001000111",  -- sqrt(5007) = 71
"001000111",  -- sqrt(5008) = 71
"001000111",  -- sqrt(5009) = 71
"001000111",  -- sqrt(5010) = 71
"001000111",  -- sqrt(5011) = 71
"001000111",  -- sqrt(5012) = 71
"001000111",  -- sqrt(5013) = 71
"001000111",  -- sqrt(5014) = 71
"001000111",  -- sqrt(5015) = 71
"001000111",  -- sqrt(5016) = 71
"001000111",  -- sqrt(5017) = 71
"001000111",  -- sqrt(5018) = 71
"001000111",  -- sqrt(5019) = 71
"001000111",  -- sqrt(5020) = 71
"001000111",  -- sqrt(5021) = 71
"001000111",  -- sqrt(5022) = 71
"001000111",  -- sqrt(5023) = 71
"001000111",  -- sqrt(5024) = 71
"001000111",  -- sqrt(5025) = 71
"001000111",  -- sqrt(5026) = 71
"001000111",  -- sqrt(5027) = 71
"001000111",  -- sqrt(5028) = 71
"001000111",  -- sqrt(5029) = 71
"001000111",  -- sqrt(5030) = 71
"001000111",  -- sqrt(5031) = 71
"001000111",  -- sqrt(5032) = 71
"001000111",  -- sqrt(5033) = 71
"001000111",  -- sqrt(5034) = 71
"001000111",  -- sqrt(5035) = 71
"001000111",  -- sqrt(5036) = 71
"001000111",  -- sqrt(5037) = 71
"001000111",  -- sqrt(5038) = 71
"001000111",  -- sqrt(5039) = 71
"001000111",  -- sqrt(5040) = 71
"001000111",  -- sqrt(5041) = 71
"001000111",  -- sqrt(5042) = 71
"001000111",  -- sqrt(5043) = 71
"001000111",  -- sqrt(5044) = 71
"001000111",  -- sqrt(5045) = 71
"001000111",  -- sqrt(5046) = 71
"001000111",  -- sqrt(5047) = 71
"001000111",  -- sqrt(5048) = 71
"001000111",  -- sqrt(5049) = 71
"001000111",  -- sqrt(5050) = 71
"001000111",  -- sqrt(5051) = 71
"001000111",  -- sqrt(5052) = 71
"001000111",  -- sqrt(5053) = 71
"001000111",  -- sqrt(5054) = 71
"001000111",  -- sqrt(5055) = 71
"001000111",  -- sqrt(5056) = 71
"001000111",  -- sqrt(5057) = 71
"001000111",  -- sqrt(5058) = 71
"001000111",  -- sqrt(5059) = 71
"001000111",  -- sqrt(5060) = 71
"001000111",  -- sqrt(5061) = 71
"001000111",  -- sqrt(5062) = 71
"001000111",  -- sqrt(5063) = 71
"001000111",  -- sqrt(5064) = 71
"001000111",  -- sqrt(5065) = 71
"001000111",  -- sqrt(5066) = 71
"001000111",  -- sqrt(5067) = 71
"001000111",  -- sqrt(5068) = 71
"001000111",  -- sqrt(5069) = 71
"001000111",  -- sqrt(5070) = 71
"001000111",  -- sqrt(5071) = 71
"001000111",  -- sqrt(5072) = 71
"001000111",  -- sqrt(5073) = 71
"001000111",  -- sqrt(5074) = 71
"001000111",  -- sqrt(5075) = 71
"001000111",  -- sqrt(5076) = 71
"001000111",  -- sqrt(5077) = 71
"001000111",  -- sqrt(5078) = 71
"001000111",  -- sqrt(5079) = 71
"001000111",  -- sqrt(5080) = 71
"001000111",  -- sqrt(5081) = 71
"001000111",  -- sqrt(5082) = 71
"001000111",  -- sqrt(5083) = 71
"001000111",  -- sqrt(5084) = 71
"001000111",  -- sqrt(5085) = 71
"001000111",  -- sqrt(5086) = 71
"001000111",  -- sqrt(5087) = 71
"001000111",  -- sqrt(5088) = 71
"001000111",  -- sqrt(5089) = 71
"001000111",  -- sqrt(5090) = 71
"001000111",  -- sqrt(5091) = 71
"001000111",  -- sqrt(5092) = 71
"001000111",  -- sqrt(5093) = 71
"001000111",  -- sqrt(5094) = 71
"001000111",  -- sqrt(5095) = 71
"001000111",  -- sqrt(5096) = 71
"001000111",  -- sqrt(5097) = 71
"001000111",  -- sqrt(5098) = 71
"001000111",  -- sqrt(5099) = 71
"001000111",  -- sqrt(5100) = 71
"001000111",  -- sqrt(5101) = 71
"001000111",  -- sqrt(5102) = 71
"001000111",  -- sqrt(5103) = 71
"001000111",  -- sqrt(5104) = 71
"001000111",  -- sqrt(5105) = 71
"001000111",  -- sqrt(5106) = 71
"001000111",  -- sqrt(5107) = 71
"001000111",  -- sqrt(5108) = 71
"001000111",  -- sqrt(5109) = 71
"001000111",  -- sqrt(5110) = 71
"001000111",  -- sqrt(5111) = 71
"001000111",  -- sqrt(5112) = 71
"001001000",  -- sqrt(5113) = 72
"001001000",  -- sqrt(5114) = 72
"001001000",  -- sqrt(5115) = 72
"001001000",  -- sqrt(5116) = 72
"001001000",  -- sqrt(5117) = 72
"001001000",  -- sqrt(5118) = 72
"001001000",  -- sqrt(5119) = 72
"001001000",  -- sqrt(5120) = 72
"001001000",  -- sqrt(5121) = 72
"001001000",  -- sqrt(5122) = 72
"001001000",  -- sqrt(5123) = 72
"001001000",  -- sqrt(5124) = 72
"001001000",  -- sqrt(5125) = 72
"001001000",  -- sqrt(5126) = 72
"001001000",  -- sqrt(5127) = 72
"001001000",  -- sqrt(5128) = 72
"001001000",  -- sqrt(5129) = 72
"001001000",  -- sqrt(5130) = 72
"001001000",  -- sqrt(5131) = 72
"001001000",  -- sqrt(5132) = 72
"001001000",  -- sqrt(5133) = 72
"001001000",  -- sqrt(5134) = 72
"001001000",  -- sqrt(5135) = 72
"001001000",  -- sqrt(5136) = 72
"001001000",  -- sqrt(5137) = 72
"001001000",  -- sqrt(5138) = 72
"001001000",  -- sqrt(5139) = 72
"001001000",  -- sqrt(5140) = 72
"001001000",  -- sqrt(5141) = 72
"001001000",  -- sqrt(5142) = 72
"001001000",  -- sqrt(5143) = 72
"001001000",  -- sqrt(5144) = 72
"001001000",  -- sqrt(5145) = 72
"001001000",  -- sqrt(5146) = 72
"001001000",  -- sqrt(5147) = 72
"001001000",  -- sqrt(5148) = 72
"001001000",  -- sqrt(5149) = 72
"001001000",  -- sqrt(5150) = 72
"001001000",  -- sqrt(5151) = 72
"001001000",  -- sqrt(5152) = 72
"001001000",  -- sqrt(5153) = 72
"001001000",  -- sqrt(5154) = 72
"001001000",  -- sqrt(5155) = 72
"001001000",  -- sqrt(5156) = 72
"001001000",  -- sqrt(5157) = 72
"001001000",  -- sqrt(5158) = 72
"001001000",  -- sqrt(5159) = 72
"001001000",  -- sqrt(5160) = 72
"001001000",  -- sqrt(5161) = 72
"001001000",  -- sqrt(5162) = 72
"001001000",  -- sqrt(5163) = 72
"001001000",  -- sqrt(5164) = 72
"001001000",  -- sqrt(5165) = 72
"001001000",  -- sqrt(5166) = 72
"001001000",  -- sqrt(5167) = 72
"001001000",  -- sqrt(5168) = 72
"001001000",  -- sqrt(5169) = 72
"001001000",  -- sqrt(5170) = 72
"001001000",  -- sqrt(5171) = 72
"001001000",  -- sqrt(5172) = 72
"001001000",  -- sqrt(5173) = 72
"001001000",  -- sqrt(5174) = 72
"001001000",  -- sqrt(5175) = 72
"001001000",  -- sqrt(5176) = 72
"001001000",  -- sqrt(5177) = 72
"001001000",  -- sqrt(5178) = 72
"001001000",  -- sqrt(5179) = 72
"001001000",  -- sqrt(5180) = 72
"001001000",  -- sqrt(5181) = 72
"001001000",  -- sqrt(5182) = 72
"001001000",  -- sqrt(5183) = 72
"001001000",  -- sqrt(5184) = 72
"001001000",  -- sqrt(5185) = 72
"001001000",  -- sqrt(5186) = 72
"001001000",  -- sqrt(5187) = 72
"001001000",  -- sqrt(5188) = 72
"001001000",  -- sqrt(5189) = 72
"001001000",  -- sqrt(5190) = 72
"001001000",  -- sqrt(5191) = 72
"001001000",  -- sqrt(5192) = 72
"001001000",  -- sqrt(5193) = 72
"001001000",  -- sqrt(5194) = 72
"001001000",  -- sqrt(5195) = 72
"001001000",  -- sqrt(5196) = 72
"001001000",  -- sqrt(5197) = 72
"001001000",  -- sqrt(5198) = 72
"001001000",  -- sqrt(5199) = 72
"001001000",  -- sqrt(5200) = 72
"001001000",  -- sqrt(5201) = 72
"001001000",  -- sqrt(5202) = 72
"001001000",  -- sqrt(5203) = 72
"001001000",  -- sqrt(5204) = 72
"001001000",  -- sqrt(5205) = 72
"001001000",  -- sqrt(5206) = 72
"001001000",  -- sqrt(5207) = 72
"001001000",  -- sqrt(5208) = 72
"001001000",  -- sqrt(5209) = 72
"001001000",  -- sqrt(5210) = 72
"001001000",  -- sqrt(5211) = 72
"001001000",  -- sqrt(5212) = 72
"001001000",  -- sqrt(5213) = 72
"001001000",  -- sqrt(5214) = 72
"001001000",  -- sqrt(5215) = 72
"001001000",  -- sqrt(5216) = 72
"001001000",  -- sqrt(5217) = 72
"001001000",  -- sqrt(5218) = 72
"001001000",  -- sqrt(5219) = 72
"001001000",  -- sqrt(5220) = 72
"001001000",  -- sqrt(5221) = 72
"001001000",  -- sqrt(5222) = 72
"001001000",  -- sqrt(5223) = 72
"001001000",  -- sqrt(5224) = 72
"001001000",  -- sqrt(5225) = 72
"001001000",  -- sqrt(5226) = 72
"001001000",  -- sqrt(5227) = 72
"001001000",  -- sqrt(5228) = 72
"001001000",  -- sqrt(5229) = 72
"001001000",  -- sqrt(5230) = 72
"001001000",  -- sqrt(5231) = 72
"001001000",  -- sqrt(5232) = 72
"001001000",  -- sqrt(5233) = 72
"001001000",  -- sqrt(5234) = 72
"001001000",  -- sqrt(5235) = 72
"001001000",  -- sqrt(5236) = 72
"001001000",  -- sqrt(5237) = 72
"001001000",  -- sqrt(5238) = 72
"001001000",  -- sqrt(5239) = 72
"001001000",  -- sqrt(5240) = 72
"001001000",  -- sqrt(5241) = 72
"001001000",  -- sqrt(5242) = 72
"001001000",  -- sqrt(5243) = 72
"001001000",  -- sqrt(5244) = 72
"001001000",  -- sqrt(5245) = 72
"001001000",  -- sqrt(5246) = 72
"001001000",  -- sqrt(5247) = 72
"001001000",  -- sqrt(5248) = 72
"001001000",  -- sqrt(5249) = 72
"001001000",  -- sqrt(5250) = 72
"001001000",  -- sqrt(5251) = 72
"001001000",  -- sqrt(5252) = 72
"001001000",  -- sqrt(5253) = 72
"001001000",  -- sqrt(5254) = 72
"001001000",  -- sqrt(5255) = 72
"001001000",  -- sqrt(5256) = 72
"001001001",  -- sqrt(5257) = 73
"001001001",  -- sqrt(5258) = 73
"001001001",  -- sqrt(5259) = 73
"001001001",  -- sqrt(5260) = 73
"001001001",  -- sqrt(5261) = 73
"001001001",  -- sqrt(5262) = 73
"001001001",  -- sqrt(5263) = 73
"001001001",  -- sqrt(5264) = 73
"001001001",  -- sqrt(5265) = 73
"001001001",  -- sqrt(5266) = 73
"001001001",  -- sqrt(5267) = 73
"001001001",  -- sqrt(5268) = 73
"001001001",  -- sqrt(5269) = 73
"001001001",  -- sqrt(5270) = 73
"001001001",  -- sqrt(5271) = 73
"001001001",  -- sqrt(5272) = 73
"001001001",  -- sqrt(5273) = 73
"001001001",  -- sqrt(5274) = 73
"001001001",  -- sqrt(5275) = 73
"001001001",  -- sqrt(5276) = 73
"001001001",  -- sqrt(5277) = 73
"001001001",  -- sqrt(5278) = 73
"001001001",  -- sqrt(5279) = 73
"001001001",  -- sqrt(5280) = 73
"001001001",  -- sqrt(5281) = 73
"001001001",  -- sqrt(5282) = 73
"001001001",  -- sqrt(5283) = 73
"001001001",  -- sqrt(5284) = 73
"001001001",  -- sqrt(5285) = 73
"001001001",  -- sqrt(5286) = 73
"001001001",  -- sqrt(5287) = 73
"001001001",  -- sqrt(5288) = 73
"001001001",  -- sqrt(5289) = 73
"001001001",  -- sqrt(5290) = 73
"001001001",  -- sqrt(5291) = 73
"001001001",  -- sqrt(5292) = 73
"001001001",  -- sqrt(5293) = 73
"001001001",  -- sqrt(5294) = 73
"001001001",  -- sqrt(5295) = 73
"001001001",  -- sqrt(5296) = 73
"001001001",  -- sqrt(5297) = 73
"001001001",  -- sqrt(5298) = 73
"001001001",  -- sqrt(5299) = 73
"001001001",  -- sqrt(5300) = 73
"001001001",  -- sqrt(5301) = 73
"001001001",  -- sqrt(5302) = 73
"001001001",  -- sqrt(5303) = 73
"001001001",  -- sqrt(5304) = 73
"001001001",  -- sqrt(5305) = 73
"001001001",  -- sqrt(5306) = 73
"001001001",  -- sqrt(5307) = 73
"001001001",  -- sqrt(5308) = 73
"001001001",  -- sqrt(5309) = 73
"001001001",  -- sqrt(5310) = 73
"001001001",  -- sqrt(5311) = 73
"001001001",  -- sqrt(5312) = 73
"001001001",  -- sqrt(5313) = 73
"001001001",  -- sqrt(5314) = 73
"001001001",  -- sqrt(5315) = 73
"001001001",  -- sqrt(5316) = 73
"001001001",  -- sqrt(5317) = 73
"001001001",  -- sqrt(5318) = 73
"001001001",  -- sqrt(5319) = 73
"001001001",  -- sqrt(5320) = 73
"001001001",  -- sqrt(5321) = 73
"001001001",  -- sqrt(5322) = 73
"001001001",  -- sqrt(5323) = 73
"001001001",  -- sqrt(5324) = 73
"001001001",  -- sqrt(5325) = 73
"001001001",  -- sqrt(5326) = 73
"001001001",  -- sqrt(5327) = 73
"001001001",  -- sqrt(5328) = 73
"001001001",  -- sqrt(5329) = 73
"001001001",  -- sqrt(5330) = 73
"001001001",  -- sqrt(5331) = 73
"001001001",  -- sqrt(5332) = 73
"001001001",  -- sqrt(5333) = 73
"001001001",  -- sqrt(5334) = 73
"001001001",  -- sqrt(5335) = 73
"001001001",  -- sqrt(5336) = 73
"001001001",  -- sqrt(5337) = 73
"001001001",  -- sqrt(5338) = 73
"001001001",  -- sqrt(5339) = 73
"001001001",  -- sqrt(5340) = 73
"001001001",  -- sqrt(5341) = 73
"001001001",  -- sqrt(5342) = 73
"001001001",  -- sqrt(5343) = 73
"001001001",  -- sqrt(5344) = 73
"001001001",  -- sqrt(5345) = 73
"001001001",  -- sqrt(5346) = 73
"001001001",  -- sqrt(5347) = 73
"001001001",  -- sqrt(5348) = 73
"001001001",  -- sqrt(5349) = 73
"001001001",  -- sqrt(5350) = 73
"001001001",  -- sqrt(5351) = 73
"001001001",  -- sqrt(5352) = 73
"001001001",  -- sqrt(5353) = 73
"001001001",  -- sqrt(5354) = 73
"001001001",  -- sqrt(5355) = 73
"001001001",  -- sqrt(5356) = 73
"001001001",  -- sqrt(5357) = 73
"001001001",  -- sqrt(5358) = 73
"001001001",  -- sqrt(5359) = 73
"001001001",  -- sqrt(5360) = 73
"001001001",  -- sqrt(5361) = 73
"001001001",  -- sqrt(5362) = 73
"001001001",  -- sqrt(5363) = 73
"001001001",  -- sqrt(5364) = 73
"001001001",  -- sqrt(5365) = 73
"001001001",  -- sqrt(5366) = 73
"001001001",  -- sqrt(5367) = 73
"001001001",  -- sqrt(5368) = 73
"001001001",  -- sqrt(5369) = 73
"001001001",  -- sqrt(5370) = 73
"001001001",  -- sqrt(5371) = 73
"001001001",  -- sqrt(5372) = 73
"001001001",  -- sqrt(5373) = 73
"001001001",  -- sqrt(5374) = 73
"001001001",  -- sqrt(5375) = 73
"001001001",  -- sqrt(5376) = 73
"001001001",  -- sqrt(5377) = 73
"001001001",  -- sqrt(5378) = 73
"001001001",  -- sqrt(5379) = 73
"001001001",  -- sqrt(5380) = 73
"001001001",  -- sqrt(5381) = 73
"001001001",  -- sqrt(5382) = 73
"001001001",  -- sqrt(5383) = 73
"001001001",  -- sqrt(5384) = 73
"001001001",  -- sqrt(5385) = 73
"001001001",  -- sqrt(5386) = 73
"001001001",  -- sqrt(5387) = 73
"001001001",  -- sqrt(5388) = 73
"001001001",  -- sqrt(5389) = 73
"001001001",  -- sqrt(5390) = 73
"001001001",  -- sqrt(5391) = 73
"001001001",  -- sqrt(5392) = 73
"001001001",  -- sqrt(5393) = 73
"001001001",  -- sqrt(5394) = 73
"001001001",  -- sqrt(5395) = 73
"001001001",  -- sqrt(5396) = 73
"001001001",  -- sqrt(5397) = 73
"001001001",  -- sqrt(5398) = 73
"001001001",  -- sqrt(5399) = 73
"001001001",  -- sqrt(5400) = 73
"001001001",  -- sqrt(5401) = 73
"001001001",  -- sqrt(5402) = 73
"001001010",  -- sqrt(5403) = 74
"001001010",  -- sqrt(5404) = 74
"001001010",  -- sqrt(5405) = 74
"001001010",  -- sqrt(5406) = 74
"001001010",  -- sqrt(5407) = 74
"001001010",  -- sqrt(5408) = 74
"001001010",  -- sqrt(5409) = 74
"001001010",  -- sqrt(5410) = 74
"001001010",  -- sqrt(5411) = 74
"001001010",  -- sqrt(5412) = 74
"001001010",  -- sqrt(5413) = 74
"001001010",  -- sqrt(5414) = 74
"001001010",  -- sqrt(5415) = 74
"001001010",  -- sqrt(5416) = 74
"001001010",  -- sqrt(5417) = 74
"001001010",  -- sqrt(5418) = 74
"001001010",  -- sqrt(5419) = 74
"001001010",  -- sqrt(5420) = 74
"001001010",  -- sqrt(5421) = 74
"001001010",  -- sqrt(5422) = 74
"001001010",  -- sqrt(5423) = 74
"001001010",  -- sqrt(5424) = 74
"001001010",  -- sqrt(5425) = 74
"001001010",  -- sqrt(5426) = 74
"001001010",  -- sqrt(5427) = 74
"001001010",  -- sqrt(5428) = 74
"001001010",  -- sqrt(5429) = 74
"001001010",  -- sqrt(5430) = 74
"001001010",  -- sqrt(5431) = 74
"001001010",  -- sqrt(5432) = 74
"001001010",  -- sqrt(5433) = 74
"001001010",  -- sqrt(5434) = 74
"001001010",  -- sqrt(5435) = 74
"001001010",  -- sqrt(5436) = 74
"001001010",  -- sqrt(5437) = 74
"001001010",  -- sqrt(5438) = 74
"001001010",  -- sqrt(5439) = 74
"001001010",  -- sqrt(5440) = 74
"001001010",  -- sqrt(5441) = 74
"001001010",  -- sqrt(5442) = 74
"001001010",  -- sqrt(5443) = 74
"001001010",  -- sqrt(5444) = 74
"001001010",  -- sqrt(5445) = 74
"001001010",  -- sqrt(5446) = 74
"001001010",  -- sqrt(5447) = 74
"001001010",  -- sqrt(5448) = 74
"001001010",  -- sqrt(5449) = 74
"001001010",  -- sqrt(5450) = 74
"001001010",  -- sqrt(5451) = 74
"001001010",  -- sqrt(5452) = 74
"001001010",  -- sqrt(5453) = 74
"001001010",  -- sqrt(5454) = 74
"001001010",  -- sqrt(5455) = 74
"001001010",  -- sqrt(5456) = 74
"001001010",  -- sqrt(5457) = 74
"001001010",  -- sqrt(5458) = 74
"001001010",  -- sqrt(5459) = 74
"001001010",  -- sqrt(5460) = 74
"001001010",  -- sqrt(5461) = 74
"001001010",  -- sqrt(5462) = 74
"001001010",  -- sqrt(5463) = 74
"001001010",  -- sqrt(5464) = 74
"001001010",  -- sqrt(5465) = 74
"001001010",  -- sqrt(5466) = 74
"001001010",  -- sqrt(5467) = 74
"001001010",  -- sqrt(5468) = 74
"001001010",  -- sqrt(5469) = 74
"001001010",  -- sqrt(5470) = 74
"001001010",  -- sqrt(5471) = 74
"001001010",  -- sqrt(5472) = 74
"001001010",  -- sqrt(5473) = 74
"001001010",  -- sqrt(5474) = 74
"001001010",  -- sqrt(5475) = 74
"001001010",  -- sqrt(5476) = 74
"001001010",  -- sqrt(5477) = 74
"001001010",  -- sqrt(5478) = 74
"001001010",  -- sqrt(5479) = 74
"001001010",  -- sqrt(5480) = 74
"001001010",  -- sqrt(5481) = 74
"001001010",  -- sqrt(5482) = 74
"001001010",  -- sqrt(5483) = 74
"001001010",  -- sqrt(5484) = 74
"001001010",  -- sqrt(5485) = 74
"001001010",  -- sqrt(5486) = 74
"001001010",  -- sqrt(5487) = 74
"001001010",  -- sqrt(5488) = 74
"001001010",  -- sqrt(5489) = 74
"001001010",  -- sqrt(5490) = 74
"001001010",  -- sqrt(5491) = 74
"001001010",  -- sqrt(5492) = 74
"001001010",  -- sqrt(5493) = 74
"001001010",  -- sqrt(5494) = 74
"001001010",  -- sqrt(5495) = 74
"001001010",  -- sqrt(5496) = 74
"001001010",  -- sqrt(5497) = 74
"001001010",  -- sqrt(5498) = 74
"001001010",  -- sqrt(5499) = 74
"001001010",  -- sqrt(5500) = 74
"001001010",  -- sqrt(5501) = 74
"001001010",  -- sqrt(5502) = 74
"001001010",  -- sqrt(5503) = 74
"001001010",  -- sqrt(5504) = 74
"001001010",  -- sqrt(5505) = 74
"001001010",  -- sqrt(5506) = 74
"001001010",  -- sqrt(5507) = 74
"001001010",  -- sqrt(5508) = 74
"001001010",  -- sqrt(5509) = 74
"001001010",  -- sqrt(5510) = 74
"001001010",  -- sqrt(5511) = 74
"001001010",  -- sqrt(5512) = 74
"001001010",  -- sqrt(5513) = 74
"001001010",  -- sqrt(5514) = 74
"001001010",  -- sqrt(5515) = 74
"001001010",  -- sqrt(5516) = 74
"001001010",  -- sqrt(5517) = 74
"001001010",  -- sqrt(5518) = 74
"001001010",  -- sqrt(5519) = 74
"001001010",  -- sqrt(5520) = 74
"001001010",  -- sqrt(5521) = 74
"001001010",  -- sqrt(5522) = 74
"001001010",  -- sqrt(5523) = 74
"001001010",  -- sqrt(5524) = 74
"001001010",  -- sqrt(5525) = 74
"001001010",  -- sqrt(5526) = 74
"001001010",  -- sqrt(5527) = 74
"001001010",  -- sqrt(5528) = 74
"001001010",  -- sqrt(5529) = 74
"001001010",  -- sqrt(5530) = 74
"001001010",  -- sqrt(5531) = 74
"001001010",  -- sqrt(5532) = 74
"001001010",  -- sqrt(5533) = 74
"001001010",  -- sqrt(5534) = 74
"001001010",  -- sqrt(5535) = 74
"001001010",  -- sqrt(5536) = 74
"001001010",  -- sqrt(5537) = 74
"001001010",  -- sqrt(5538) = 74
"001001010",  -- sqrt(5539) = 74
"001001010",  -- sqrt(5540) = 74
"001001010",  -- sqrt(5541) = 74
"001001010",  -- sqrt(5542) = 74
"001001010",  -- sqrt(5543) = 74
"001001010",  -- sqrt(5544) = 74
"001001010",  -- sqrt(5545) = 74
"001001010",  -- sqrt(5546) = 74
"001001010",  -- sqrt(5547) = 74
"001001010",  -- sqrt(5548) = 74
"001001010",  -- sqrt(5549) = 74
"001001010",  -- sqrt(5550) = 74
"001001011",  -- sqrt(5551) = 75
"001001011",  -- sqrt(5552) = 75
"001001011",  -- sqrt(5553) = 75
"001001011",  -- sqrt(5554) = 75
"001001011",  -- sqrt(5555) = 75
"001001011",  -- sqrt(5556) = 75
"001001011",  -- sqrt(5557) = 75
"001001011",  -- sqrt(5558) = 75
"001001011",  -- sqrt(5559) = 75
"001001011",  -- sqrt(5560) = 75
"001001011",  -- sqrt(5561) = 75
"001001011",  -- sqrt(5562) = 75
"001001011",  -- sqrt(5563) = 75
"001001011",  -- sqrt(5564) = 75
"001001011",  -- sqrt(5565) = 75
"001001011",  -- sqrt(5566) = 75
"001001011",  -- sqrt(5567) = 75
"001001011",  -- sqrt(5568) = 75
"001001011",  -- sqrt(5569) = 75
"001001011",  -- sqrt(5570) = 75
"001001011",  -- sqrt(5571) = 75
"001001011",  -- sqrt(5572) = 75
"001001011",  -- sqrt(5573) = 75
"001001011",  -- sqrt(5574) = 75
"001001011",  -- sqrt(5575) = 75
"001001011",  -- sqrt(5576) = 75
"001001011",  -- sqrt(5577) = 75
"001001011",  -- sqrt(5578) = 75
"001001011",  -- sqrt(5579) = 75
"001001011",  -- sqrt(5580) = 75
"001001011",  -- sqrt(5581) = 75
"001001011",  -- sqrt(5582) = 75
"001001011",  -- sqrt(5583) = 75
"001001011",  -- sqrt(5584) = 75
"001001011",  -- sqrt(5585) = 75
"001001011",  -- sqrt(5586) = 75
"001001011",  -- sqrt(5587) = 75
"001001011",  -- sqrt(5588) = 75
"001001011",  -- sqrt(5589) = 75
"001001011",  -- sqrt(5590) = 75
"001001011",  -- sqrt(5591) = 75
"001001011",  -- sqrt(5592) = 75
"001001011",  -- sqrt(5593) = 75
"001001011",  -- sqrt(5594) = 75
"001001011",  -- sqrt(5595) = 75
"001001011",  -- sqrt(5596) = 75
"001001011",  -- sqrt(5597) = 75
"001001011",  -- sqrt(5598) = 75
"001001011",  -- sqrt(5599) = 75
"001001011",  -- sqrt(5600) = 75
"001001011",  -- sqrt(5601) = 75
"001001011",  -- sqrt(5602) = 75
"001001011",  -- sqrt(5603) = 75
"001001011",  -- sqrt(5604) = 75
"001001011",  -- sqrt(5605) = 75
"001001011",  -- sqrt(5606) = 75
"001001011",  -- sqrt(5607) = 75
"001001011",  -- sqrt(5608) = 75
"001001011",  -- sqrt(5609) = 75
"001001011",  -- sqrt(5610) = 75
"001001011",  -- sqrt(5611) = 75
"001001011",  -- sqrt(5612) = 75
"001001011",  -- sqrt(5613) = 75
"001001011",  -- sqrt(5614) = 75
"001001011",  -- sqrt(5615) = 75
"001001011",  -- sqrt(5616) = 75
"001001011",  -- sqrt(5617) = 75
"001001011",  -- sqrt(5618) = 75
"001001011",  -- sqrt(5619) = 75
"001001011",  -- sqrt(5620) = 75
"001001011",  -- sqrt(5621) = 75
"001001011",  -- sqrt(5622) = 75
"001001011",  -- sqrt(5623) = 75
"001001011",  -- sqrt(5624) = 75
"001001011",  -- sqrt(5625) = 75
"001001011",  -- sqrt(5626) = 75
"001001011",  -- sqrt(5627) = 75
"001001011",  -- sqrt(5628) = 75
"001001011",  -- sqrt(5629) = 75
"001001011",  -- sqrt(5630) = 75
"001001011",  -- sqrt(5631) = 75
"001001011",  -- sqrt(5632) = 75
"001001011",  -- sqrt(5633) = 75
"001001011",  -- sqrt(5634) = 75
"001001011",  -- sqrt(5635) = 75
"001001011",  -- sqrt(5636) = 75
"001001011",  -- sqrt(5637) = 75
"001001011",  -- sqrt(5638) = 75
"001001011",  -- sqrt(5639) = 75
"001001011",  -- sqrt(5640) = 75
"001001011",  -- sqrt(5641) = 75
"001001011",  -- sqrt(5642) = 75
"001001011",  -- sqrt(5643) = 75
"001001011",  -- sqrt(5644) = 75
"001001011",  -- sqrt(5645) = 75
"001001011",  -- sqrt(5646) = 75
"001001011",  -- sqrt(5647) = 75
"001001011",  -- sqrt(5648) = 75
"001001011",  -- sqrt(5649) = 75
"001001011",  -- sqrt(5650) = 75
"001001011",  -- sqrt(5651) = 75
"001001011",  -- sqrt(5652) = 75
"001001011",  -- sqrt(5653) = 75
"001001011",  -- sqrt(5654) = 75
"001001011",  -- sqrt(5655) = 75
"001001011",  -- sqrt(5656) = 75
"001001011",  -- sqrt(5657) = 75
"001001011",  -- sqrt(5658) = 75
"001001011",  -- sqrt(5659) = 75
"001001011",  -- sqrt(5660) = 75
"001001011",  -- sqrt(5661) = 75
"001001011",  -- sqrt(5662) = 75
"001001011",  -- sqrt(5663) = 75
"001001011",  -- sqrt(5664) = 75
"001001011",  -- sqrt(5665) = 75
"001001011",  -- sqrt(5666) = 75
"001001011",  -- sqrt(5667) = 75
"001001011",  -- sqrt(5668) = 75
"001001011",  -- sqrt(5669) = 75
"001001011",  -- sqrt(5670) = 75
"001001011",  -- sqrt(5671) = 75
"001001011",  -- sqrt(5672) = 75
"001001011",  -- sqrt(5673) = 75
"001001011",  -- sqrt(5674) = 75
"001001011",  -- sqrt(5675) = 75
"001001011",  -- sqrt(5676) = 75
"001001011",  -- sqrt(5677) = 75
"001001011",  -- sqrt(5678) = 75
"001001011",  -- sqrt(5679) = 75
"001001011",  -- sqrt(5680) = 75
"001001011",  -- sqrt(5681) = 75
"001001011",  -- sqrt(5682) = 75
"001001011",  -- sqrt(5683) = 75
"001001011",  -- sqrt(5684) = 75
"001001011",  -- sqrt(5685) = 75
"001001011",  -- sqrt(5686) = 75
"001001011",  -- sqrt(5687) = 75
"001001011",  -- sqrt(5688) = 75
"001001011",  -- sqrt(5689) = 75
"001001011",  -- sqrt(5690) = 75
"001001011",  -- sqrt(5691) = 75
"001001011",  -- sqrt(5692) = 75
"001001011",  -- sqrt(5693) = 75
"001001011",  -- sqrt(5694) = 75
"001001011",  -- sqrt(5695) = 75
"001001011",  -- sqrt(5696) = 75
"001001011",  -- sqrt(5697) = 75
"001001011",  -- sqrt(5698) = 75
"001001011",  -- sqrt(5699) = 75
"001001011",  -- sqrt(5700) = 75
"001001100",  -- sqrt(5701) = 76
"001001100",  -- sqrt(5702) = 76
"001001100",  -- sqrt(5703) = 76
"001001100",  -- sqrt(5704) = 76
"001001100",  -- sqrt(5705) = 76
"001001100",  -- sqrt(5706) = 76
"001001100",  -- sqrt(5707) = 76
"001001100",  -- sqrt(5708) = 76
"001001100",  -- sqrt(5709) = 76
"001001100",  -- sqrt(5710) = 76
"001001100",  -- sqrt(5711) = 76
"001001100",  -- sqrt(5712) = 76
"001001100",  -- sqrt(5713) = 76
"001001100",  -- sqrt(5714) = 76
"001001100",  -- sqrt(5715) = 76
"001001100",  -- sqrt(5716) = 76
"001001100",  -- sqrt(5717) = 76
"001001100",  -- sqrt(5718) = 76
"001001100",  -- sqrt(5719) = 76
"001001100",  -- sqrt(5720) = 76
"001001100",  -- sqrt(5721) = 76
"001001100",  -- sqrt(5722) = 76
"001001100",  -- sqrt(5723) = 76
"001001100",  -- sqrt(5724) = 76
"001001100",  -- sqrt(5725) = 76
"001001100",  -- sqrt(5726) = 76
"001001100",  -- sqrt(5727) = 76
"001001100",  -- sqrt(5728) = 76
"001001100",  -- sqrt(5729) = 76
"001001100",  -- sqrt(5730) = 76
"001001100",  -- sqrt(5731) = 76
"001001100",  -- sqrt(5732) = 76
"001001100",  -- sqrt(5733) = 76
"001001100",  -- sqrt(5734) = 76
"001001100",  -- sqrt(5735) = 76
"001001100",  -- sqrt(5736) = 76
"001001100",  -- sqrt(5737) = 76
"001001100",  -- sqrt(5738) = 76
"001001100",  -- sqrt(5739) = 76
"001001100",  -- sqrt(5740) = 76
"001001100",  -- sqrt(5741) = 76
"001001100",  -- sqrt(5742) = 76
"001001100",  -- sqrt(5743) = 76
"001001100",  -- sqrt(5744) = 76
"001001100",  -- sqrt(5745) = 76
"001001100",  -- sqrt(5746) = 76
"001001100",  -- sqrt(5747) = 76
"001001100",  -- sqrt(5748) = 76
"001001100",  -- sqrt(5749) = 76
"001001100",  -- sqrt(5750) = 76
"001001100",  -- sqrt(5751) = 76
"001001100",  -- sqrt(5752) = 76
"001001100",  -- sqrt(5753) = 76
"001001100",  -- sqrt(5754) = 76
"001001100",  -- sqrt(5755) = 76
"001001100",  -- sqrt(5756) = 76
"001001100",  -- sqrt(5757) = 76
"001001100",  -- sqrt(5758) = 76
"001001100",  -- sqrt(5759) = 76
"001001100",  -- sqrt(5760) = 76
"001001100",  -- sqrt(5761) = 76
"001001100",  -- sqrt(5762) = 76
"001001100",  -- sqrt(5763) = 76
"001001100",  -- sqrt(5764) = 76
"001001100",  -- sqrt(5765) = 76
"001001100",  -- sqrt(5766) = 76
"001001100",  -- sqrt(5767) = 76
"001001100",  -- sqrt(5768) = 76
"001001100",  -- sqrt(5769) = 76
"001001100",  -- sqrt(5770) = 76
"001001100",  -- sqrt(5771) = 76
"001001100",  -- sqrt(5772) = 76
"001001100",  -- sqrt(5773) = 76
"001001100",  -- sqrt(5774) = 76
"001001100",  -- sqrt(5775) = 76
"001001100",  -- sqrt(5776) = 76
"001001100",  -- sqrt(5777) = 76
"001001100",  -- sqrt(5778) = 76
"001001100",  -- sqrt(5779) = 76
"001001100",  -- sqrt(5780) = 76
"001001100",  -- sqrt(5781) = 76
"001001100",  -- sqrt(5782) = 76
"001001100",  -- sqrt(5783) = 76
"001001100",  -- sqrt(5784) = 76
"001001100",  -- sqrt(5785) = 76
"001001100",  -- sqrt(5786) = 76
"001001100",  -- sqrt(5787) = 76
"001001100",  -- sqrt(5788) = 76
"001001100",  -- sqrt(5789) = 76
"001001100",  -- sqrt(5790) = 76
"001001100",  -- sqrt(5791) = 76
"001001100",  -- sqrt(5792) = 76
"001001100",  -- sqrt(5793) = 76
"001001100",  -- sqrt(5794) = 76
"001001100",  -- sqrt(5795) = 76
"001001100",  -- sqrt(5796) = 76
"001001100",  -- sqrt(5797) = 76
"001001100",  -- sqrt(5798) = 76
"001001100",  -- sqrt(5799) = 76
"001001100",  -- sqrt(5800) = 76
"001001100",  -- sqrt(5801) = 76
"001001100",  -- sqrt(5802) = 76
"001001100",  -- sqrt(5803) = 76
"001001100",  -- sqrt(5804) = 76
"001001100",  -- sqrt(5805) = 76
"001001100",  -- sqrt(5806) = 76
"001001100",  -- sqrt(5807) = 76
"001001100",  -- sqrt(5808) = 76
"001001100",  -- sqrt(5809) = 76
"001001100",  -- sqrt(5810) = 76
"001001100",  -- sqrt(5811) = 76
"001001100",  -- sqrt(5812) = 76
"001001100",  -- sqrt(5813) = 76
"001001100",  -- sqrt(5814) = 76
"001001100",  -- sqrt(5815) = 76
"001001100",  -- sqrt(5816) = 76
"001001100",  -- sqrt(5817) = 76
"001001100",  -- sqrt(5818) = 76
"001001100",  -- sqrt(5819) = 76
"001001100",  -- sqrt(5820) = 76
"001001100",  -- sqrt(5821) = 76
"001001100",  -- sqrt(5822) = 76
"001001100",  -- sqrt(5823) = 76
"001001100",  -- sqrt(5824) = 76
"001001100",  -- sqrt(5825) = 76
"001001100",  -- sqrt(5826) = 76
"001001100",  -- sqrt(5827) = 76
"001001100",  -- sqrt(5828) = 76
"001001100",  -- sqrt(5829) = 76
"001001100",  -- sqrt(5830) = 76
"001001100",  -- sqrt(5831) = 76
"001001100",  -- sqrt(5832) = 76
"001001100",  -- sqrt(5833) = 76
"001001100",  -- sqrt(5834) = 76
"001001100",  -- sqrt(5835) = 76
"001001100",  -- sqrt(5836) = 76
"001001100",  -- sqrt(5837) = 76
"001001100",  -- sqrt(5838) = 76
"001001100",  -- sqrt(5839) = 76
"001001100",  -- sqrt(5840) = 76
"001001100",  -- sqrt(5841) = 76
"001001100",  -- sqrt(5842) = 76
"001001100",  -- sqrt(5843) = 76
"001001100",  -- sqrt(5844) = 76
"001001100",  -- sqrt(5845) = 76
"001001100",  -- sqrt(5846) = 76
"001001100",  -- sqrt(5847) = 76
"001001100",  -- sqrt(5848) = 76
"001001100",  -- sqrt(5849) = 76
"001001100",  -- sqrt(5850) = 76
"001001100",  -- sqrt(5851) = 76
"001001100",  -- sqrt(5852) = 76
"001001101",  -- sqrt(5853) = 77
"001001101",  -- sqrt(5854) = 77
"001001101",  -- sqrt(5855) = 77
"001001101",  -- sqrt(5856) = 77
"001001101",  -- sqrt(5857) = 77
"001001101",  -- sqrt(5858) = 77
"001001101",  -- sqrt(5859) = 77
"001001101",  -- sqrt(5860) = 77
"001001101",  -- sqrt(5861) = 77
"001001101",  -- sqrt(5862) = 77
"001001101",  -- sqrt(5863) = 77
"001001101",  -- sqrt(5864) = 77
"001001101",  -- sqrt(5865) = 77
"001001101",  -- sqrt(5866) = 77
"001001101",  -- sqrt(5867) = 77
"001001101",  -- sqrt(5868) = 77
"001001101",  -- sqrt(5869) = 77
"001001101",  -- sqrt(5870) = 77
"001001101",  -- sqrt(5871) = 77
"001001101",  -- sqrt(5872) = 77
"001001101",  -- sqrt(5873) = 77
"001001101",  -- sqrt(5874) = 77
"001001101",  -- sqrt(5875) = 77
"001001101",  -- sqrt(5876) = 77
"001001101",  -- sqrt(5877) = 77
"001001101",  -- sqrt(5878) = 77
"001001101",  -- sqrt(5879) = 77
"001001101",  -- sqrt(5880) = 77
"001001101",  -- sqrt(5881) = 77
"001001101",  -- sqrt(5882) = 77
"001001101",  -- sqrt(5883) = 77
"001001101",  -- sqrt(5884) = 77
"001001101",  -- sqrt(5885) = 77
"001001101",  -- sqrt(5886) = 77
"001001101",  -- sqrt(5887) = 77
"001001101",  -- sqrt(5888) = 77
"001001101",  -- sqrt(5889) = 77
"001001101",  -- sqrt(5890) = 77
"001001101",  -- sqrt(5891) = 77
"001001101",  -- sqrt(5892) = 77
"001001101",  -- sqrt(5893) = 77
"001001101",  -- sqrt(5894) = 77
"001001101",  -- sqrt(5895) = 77
"001001101",  -- sqrt(5896) = 77
"001001101",  -- sqrt(5897) = 77
"001001101",  -- sqrt(5898) = 77
"001001101",  -- sqrt(5899) = 77
"001001101",  -- sqrt(5900) = 77
"001001101",  -- sqrt(5901) = 77
"001001101",  -- sqrt(5902) = 77
"001001101",  -- sqrt(5903) = 77
"001001101",  -- sqrt(5904) = 77
"001001101",  -- sqrt(5905) = 77
"001001101",  -- sqrt(5906) = 77
"001001101",  -- sqrt(5907) = 77
"001001101",  -- sqrt(5908) = 77
"001001101",  -- sqrt(5909) = 77
"001001101",  -- sqrt(5910) = 77
"001001101",  -- sqrt(5911) = 77
"001001101",  -- sqrt(5912) = 77
"001001101",  -- sqrt(5913) = 77
"001001101",  -- sqrt(5914) = 77
"001001101",  -- sqrt(5915) = 77
"001001101",  -- sqrt(5916) = 77
"001001101",  -- sqrt(5917) = 77
"001001101",  -- sqrt(5918) = 77
"001001101",  -- sqrt(5919) = 77
"001001101",  -- sqrt(5920) = 77
"001001101",  -- sqrt(5921) = 77
"001001101",  -- sqrt(5922) = 77
"001001101",  -- sqrt(5923) = 77
"001001101",  -- sqrt(5924) = 77
"001001101",  -- sqrt(5925) = 77
"001001101",  -- sqrt(5926) = 77
"001001101",  -- sqrt(5927) = 77
"001001101",  -- sqrt(5928) = 77
"001001101",  -- sqrt(5929) = 77
"001001101",  -- sqrt(5930) = 77
"001001101",  -- sqrt(5931) = 77
"001001101",  -- sqrt(5932) = 77
"001001101",  -- sqrt(5933) = 77
"001001101",  -- sqrt(5934) = 77
"001001101",  -- sqrt(5935) = 77
"001001101",  -- sqrt(5936) = 77
"001001101",  -- sqrt(5937) = 77
"001001101",  -- sqrt(5938) = 77
"001001101",  -- sqrt(5939) = 77
"001001101",  -- sqrt(5940) = 77
"001001101",  -- sqrt(5941) = 77
"001001101",  -- sqrt(5942) = 77
"001001101",  -- sqrt(5943) = 77
"001001101",  -- sqrt(5944) = 77
"001001101",  -- sqrt(5945) = 77
"001001101",  -- sqrt(5946) = 77
"001001101",  -- sqrt(5947) = 77
"001001101",  -- sqrt(5948) = 77
"001001101",  -- sqrt(5949) = 77
"001001101",  -- sqrt(5950) = 77
"001001101",  -- sqrt(5951) = 77
"001001101",  -- sqrt(5952) = 77
"001001101",  -- sqrt(5953) = 77
"001001101",  -- sqrt(5954) = 77
"001001101",  -- sqrt(5955) = 77
"001001101",  -- sqrt(5956) = 77
"001001101",  -- sqrt(5957) = 77
"001001101",  -- sqrt(5958) = 77
"001001101",  -- sqrt(5959) = 77
"001001101",  -- sqrt(5960) = 77
"001001101",  -- sqrt(5961) = 77
"001001101",  -- sqrt(5962) = 77
"001001101",  -- sqrt(5963) = 77
"001001101",  -- sqrt(5964) = 77
"001001101",  -- sqrt(5965) = 77
"001001101",  -- sqrt(5966) = 77
"001001101",  -- sqrt(5967) = 77
"001001101",  -- sqrt(5968) = 77
"001001101",  -- sqrt(5969) = 77
"001001101",  -- sqrt(5970) = 77
"001001101",  -- sqrt(5971) = 77
"001001101",  -- sqrt(5972) = 77
"001001101",  -- sqrt(5973) = 77
"001001101",  -- sqrt(5974) = 77
"001001101",  -- sqrt(5975) = 77
"001001101",  -- sqrt(5976) = 77
"001001101",  -- sqrt(5977) = 77
"001001101",  -- sqrt(5978) = 77
"001001101",  -- sqrt(5979) = 77
"001001101",  -- sqrt(5980) = 77
"001001101",  -- sqrt(5981) = 77
"001001101",  -- sqrt(5982) = 77
"001001101",  -- sqrt(5983) = 77
"001001101",  -- sqrt(5984) = 77
"001001101",  -- sqrt(5985) = 77
"001001101",  -- sqrt(5986) = 77
"001001101",  -- sqrt(5987) = 77
"001001101",  -- sqrt(5988) = 77
"001001101",  -- sqrt(5989) = 77
"001001101",  -- sqrt(5990) = 77
"001001101",  -- sqrt(5991) = 77
"001001101",  -- sqrt(5992) = 77
"001001101",  -- sqrt(5993) = 77
"001001101",  -- sqrt(5994) = 77
"001001101",  -- sqrt(5995) = 77
"001001101",  -- sqrt(5996) = 77
"001001101",  -- sqrt(5997) = 77
"001001101",  -- sqrt(5998) = 77
"001001101",  -- sqrt(5999) = 77
"001001101",  -- sqrt(6000) = 77
"001001101",  -- sqrt(6001) = 77
"001001101",  -- sqrt(6002) = 77
"001001101",  -- sqrt(6003) = 77
"001001101",  -- sqrt(6004) = 77
"001001101",  -- sqrt(6005) = 77
"001001101",  -- sqrt(6006) = 77
"001001110",  -- sqrt(6007) = 78
"001001110",  -- sqrt(6008) = 78
"001001110",  -- sqrt(6009) = 78
"001001110",  -- sqrt(6010) = 78
"001001110",  -- sqrt(6011) = 78
"001001110",  -- sqrt(6012) = 78
"001001110",  -- sqrt(6013) = 78
"001001110",  -- sqrt(6014) = 78
"001001110",  -- sqrt(6015) = 78
"001001110",  -- sqrt(6016) = 78
"001001110",  -- sqrt(6017) = 78
"001001110",  -- sqrt(6018) = 78
"001001110",  -- sqrt(6019) = 78
"001001110",  -- sqrt(6020) = 78
"001001110",  -- sqrt(6021) = 78
"001001110",  -- sqrt(6022) = 78
"001001110",  -- sqrt(6023) = 78
"001001110",  -- sqrt(6024) = 78
"001001110",  -- sqrt(6025) = 78
"001001110",  -- sqrt(6026) = 78
"001001110",  -- sqrt(6027) = 78
"001001110",  -- sqrt(6028) = 78
"001001110",  -- sqrt(6029) = 78
"001001110",  -- sqrt(6030) = 78
"001001110",  -- sqrt(6031) = 78
"001001110",  -- sqrt(6032) = 78
"001001110",  -- sqrt(6033) = 78
"001001110",  -- sqrt(6034) = 78
"001001110",  -- sqrt(6035) = 78
"001001110",  -- sqrt(6036) = 78
"001001110",  -- sqrt(6037) = 78
"001001110",  -- sqrt(6038) = 78
"001001110",  -- sqrt(6039) = 78
"001001110",  -- sqrt(6040) = 78
"001001110",  -- sqrt(6041) = 78
"001001110",  -- sqrt(6042) = 78
"001001110",  -- sqrt(6043) = 78
"001001110",  -- sqrt(6044) = 78
"001001110",  -- sqrt(6045) = 78
"001001110",  -- sqrt(6046) = 78
"001001110",  -- sqrt(6047) = 78
"001001110",  -- sqrt(6048) = 78
"001001110",  -- sqrt(6049) = 78
"001001110",  -- sqrt(6050) = 78
"001001110",  -- sqrt(6051) = 78
"001001110",  -- sqrt(6052) = 78
"001001110",  -- sqrt(6053) = 78
"001001110",  -- sqrt(6054) = 78
"001001110",  -- sqrt(6055) = 78
"001001110",  -- sqrt(6056) = 78
"001001110",  -- sqrt(6057) = 78
"001001110",  -- sqrt(6058) = 78
"001001110",  -- sqrt(6059) = 78
"001001110",  -- sqrt(6060) = 78
"001001110",  -- sqrt(6061) = 78
"001001110",  -- sqrt(6062) = 78
"001001110",  -- sqrt(6063) = 78
"001001110",  -- sqrt(6064) = 78
"001001110",  -- sqrt(6065) = 78
"001001110",  -- sqrt(6066) = 78
"001001110",  -- sqrt(6067) = 78
"001001110",  -- sqrt(6068) = 78
"001001110",  -- sqrt(6069) = 78
"001001110",  -- sqrt(6070) = 78
"001001110",  -- sqrt(6071) = 78
"001001110",  -- sqrt(6072) = 78
"001001110",  -- sqrt(6073) = 78
"001001110",  -- sqrt(6074) = 78
"001001110",  -- sqrt(6075) = 78
"001001110",  -- sqrt(6076) = 78
"001001110",  -- sqrt(6077) = 78
"001001110",  -- sqrt(6078) = 78
"001001110",  -- sqrt(6079) = 78
"001001110",  -- sqrt(6080) = 78
"001001110",  -- sqrt(6081) = 78
"001001110",  -- sqrt(6082) = 78
"001001110",  -- sqrt(6083) = 78
"001001110",  -- sqrt(6084) = 78
"001001110",  -- sqrt(6085) = 78
"001001110",  -- sqrt(6086) = 78
"001001110",  -- sqrt(6087) = 78
"001001110",  -- sqrt(6088) = 78
"001001110",  -- sqrt(6089) = 78
"001001110",  -- sqrt(6090) = 78
"001001110",  -- sqrt(6091) = 78
"001001110",  -- sqrt(6092) = 78
"001001110",  -- sqrt(6093) = 78
"001001110",  -- sqrt(6094) = 78
"001001110",  -- sqrt(6095) = 78
"001001110",  -- sqrt(6096) = 78
"001001110",  -- sqrt(6097) = 78
"001001110",  -- sqrt(6098) = 78
"001001110",  -- sqrt(6099) = 78
"001001110",  -- sqrt(6100) = 78
"001001110",  -- sqrt(6101) = 78
"001001110",  -- sqrt(6102) = 78
"001001110",  -- sqrt(6103) = 78
"001001110",  -- sqrt(6104) = 78
"001001110",  -- sqrt(6105) = 78
"001001110",  -- sqrt(6106) = 78
"001001110",  -- sqrt(6107) = 78
"001001110",  -- sqrt(6108) = 78
"001001110",  -- sqrt(6109) = 78
"001001110",  -- sqrt(6110) = 78
"001001110",  -- sqrt(6111) = 78
"001001110",  -- sqrt(6112) = 78
"001001110",  -- sqrt(6113) = 78
"001001110",  -- sqrt(6114) = 78
"001001110",  -- sqrt(6115) = 78
"001001110",  -- sqrt(6116) = 78
"001001110",  -- sqrt(6117) = 78
"001001110",  -- sqrt(6118) = 78
"001001110",  -- sqrt(6119) = 78
"001001110",  -- sqrt(6120) = 78
"001001110",  -- sqrt(6121) = 78
"001001110",  -- sqrt(6122) = 78
"001001110",  -- sqrt(6123) = 78
"001001110",  -- sqrt(6124) = 78
"001001110",  -- sqrt(6125) = 78
"001001110",  -- sqrt(6126) = 78
"001001110",  -- sqrt(6127) = 78
"001001110",  -- sqrt(6128) = 78
"001001110",  -- sqrt(6129) = 78
"001001110",  -- sqrt(6130) = 78
"001001110",  -- sqrt(6131) = 78
"001001110",  -- sqrt(6132) = 78
"001001110",  -- sqrt(6133) = 78
"001001110",  -- sqrt(6134) = 78
"001001110",  -- sqrt(6135) = 78
"001001110",  -- sqrt(6136) = 78
"001001110",  -- sqrt(6137) = 78
"001001110",  -- sqrt(6138) = 78
"001001110",  -- sqrt(6139) = 78
"001001110",  -- sqrt(6140) = 78
"001001110",  -- sqrt(6141) = 78
"001001110",  -- sqrt(6142) = 78
"001001110",  -- sqrt(6143) = 78
"001001110",  -- sqrt(6144) = 78
"001001110",  -- sqrt(6145) = 78
"001001110",  -- sqrt(6146) = 78
"001001110",  -- sqrt(6147) = 78
"001001110",  -- sqrt(6148) = 78
"001001110",  -- sqrt(6149) = 78
"001001110",  -- sqrt(6150) = 78
"001001110",  -- sqrt(6151) = 78
"001001110",  -- sqrt(6152) = 78
"001001110",  -- sqrt(6153) = 78
"001001110",  -- sqrt(6154) = 78
"001001110",  -- sqrt(6155) = 78
"001001110",  -- sqrt(6156) = 78
"001001110",  -- sqrt(6157) = 78
"001001110",  -- sqrt(6158) = 78
"001001110",  -- sqrt(6159) = 78
"001001110",  -- sqrt(6160) = 78
"001001110",  -- sqrt(6161) = 78
"001001110",  -- sqrt(6162) = 78
"001001111",  -- sqrt(6163) = 79
"001001111",  -- sqrt(6164) = 79
"001001111",  -- sqrt(6165) = 79
"001001111",  -- sqrt(6166) = 79
"001001111",  -- sqrt(6167) = 79
"001001111",  -- sqrt(6168) = 79
"001001111",  -- sqrt(6169) = 79
"001001111",  -- sqrt(6170) = 79
"001001111",  -- sqrt(6171) = 79
"001001111",  -- sqrt(6172) = 79
"001001111",  -- sqrt(6173) = 79
"001001111",  -- sqrt(6174) = 79
"001001111",  -- sqrt(6175) = 79
"001001111",  -- sqrt(6176) = 79
"001001111",  -- sqrt(6177) = 79
"001001111",  -- sqrt(6178) = 79
"001001111",  -- sqrt(6179) = 79
"001001111",  -- sqrt(6180) = 79
"001001111",  -- sqrt(6181) = 79
"001001111",  -- sqrt(6182) = 79
"001001111",  -- sqrt(6183) = 79
"001001111",  -- sqrt(6184) = 79
"001001111",  -- sqrt(6185) = 79
"001001111",  -- sqrt(6186) = 79
"001001111",  -- sqrt(6187) = 79
"001001111",  -- sqrt(6188) = 79
"001001111",  -- sqrt(6189) = 79
"001001111",  -- sqrt(6190) = 79
"001001111",  -- sqrt(6191) = 79
"001001111",  -- sqrt(6192) = 79
"001001111",  -- sqrt(6193) = 79
"001001111",  -- sqrt(6194) = 79
"001001111",  -- sqrt(6195) = 79
"001001111",  -- sqrt(6196) = 79
"001001111",  -- sqrt(6197) = 79
"001001111",  -- sqrt(6198) = 79
"001001111",  -- sqrt(6199) = 79
"001001111",  -- sqrt(6200) = 79
"001001111",  -- sqrt(6201) = 79
"001001111",  -- sqrt(6202) = 79
"001001111",  -- sqrt(6203) = 79
"001001111",  -- sqrt(6204) = 79
"001001111",  -- sqrt(6205) = 79
"001001111",  -- sqrt(6206) = 79
"001001111",  -- sqrt(6207) = 79
"001001111",  -- sqrt(6208) = 79
"001001111",  -- sqrt(6209) = 79
"001001111",  -- sqrt(6210) = 79
"001001111",  -- sqrt(6211) = 79
"001001111",  -- sqrt(6212) = 79
"001001111",  -- sqrt(6213) = 79
"001001111",  -- sqrt(6214) = 79
"001001111",  -- sqrt(6215) = 79
"001001111",  -- sqrt(6216) = 79
"001001111",  -- sqrt(6217) = 79
"001001111",  -- sqrt(6218) = 79
"001001111",  -- sqrt(6219) = 79
"001001111",  -- sqrt(6220) = 79
"001001111",  -- sqrt(6221) = 79
"001001111",  -- sqrt(6222) = 79
"001001111",  -- sqrt(6223) = 79
"001001111",  -- sqrt(6224) = 79
"001001111",  -- sqrt(6225) = 79
"001001111",  -- sqrt(6226) = 79
"001001111",  -- sqrt(6227) = 79
"001001111",  -- sqrt(6228) = 79
"001001111",  -- sqrt(6229) = 79
"001001111",  -- sqrt(6230) = 79
"001001111",  -- sqrt(6231) = 79
"001001111",  -- sqrt(6232) = 79
"001001111",  -- sqrt(6233) = 79
"001001111",  -- sqrt(6234) = 79
"001001111",  -- sqrt(6235) = 79
"001001111",  -- sqrt(6236) = 79
"001001111",  -- sqrt(6237) = 79
"001001111",  -- sqrt(6238) = 79
"001001111",  -- sqrt(6239) = 79
"001001111",  -- sqrt(6240) = 79
"001001111",  -- sqrt(6241) = 79
"001001111",  -- sqrt(6242) = 79
"001001111",  -- sqrt(6243) = 79
"001001111",  -- sqrt(6244) = 79
"001001111",  -- sqrt(6245) = 79
"001001111",  -- sqrt(6246) = 79
"001001111",  -- sqrt(6247) = 79
"001001111",  -- sqrt(6248) = 79
"001001111",  -- sqrt(6249) = 79
"001001111",  -- sqrt(6250) = 79
"001001111",  -- sqrt(6251) = 79
"001001111",  -- sqrt(6252) = 79
"001001111",  -- sqrt(6253) = 79
"001001111",  -- sqrt(6254) = 79
"001001111",  -- sqrt(6255) = 79
"001001111",  -- sqrt(6256) = 79
"001001111",  -- sqrt(6257) = 79
"001001111",  -- sqrt(6258) = 79
"001001111",  -- sqrt(6259) = 79
"001001111",  -- sqrt(6260) = 79
"001001111",  -- sqrt(6261) = 79
"001001111",  -- sqrt(6262) = 79
"001001111",  -- sqrt(6263) = 79
"001001111",  -- sqrt(6264) = 79
"001001111",  -- sqrt(6265) = 79
"001001111",  -- sqrt(6266) = 79
"001001111",  -- sqrt(6267) = 79
"001001111",  -- sqrt(6268) = 79
"001001111",  -- sqrt(6269) = 79
"001001111",  -- sqrt(6270) = 79
"001001111",  -- sqrt(6271) = 79
"001001111",  -- sqrt(6272) = 79
"001001111",  -- sqrt(6273) = 79
"001001111",  -- sqrt(6274) = 79
"001001111",  -- sqrt(6275) = 79
"001001111",  -- sqrt(6276) = 79
"001001111",  -- sqrt(6277) = 79
"001001111",  -- sqrt(6278) = 79
"001001111",  -- sqrt(6279) = 79
"001001111",  -- sqrt(6280) = 79
"001001111",  -- sqrt(6281) = 79
"001001111",  -- sqrt(6282) = 79
"001001111",  -- sqrt(6283) = 79
"001001111",  -- sqrt(6284) = 79
"001001111",  -- sqrt(6285) = 79
"001001111",  -- sqrt(6286) = 79
"001001111",  -- sqrt(6287) = 79
"001001111",  -- sqrt(6288) = 79
"001001111",  -- sqrt(6289) = 79
"001001111",  -- sqrt(6290) = 79
"001001111",  -- sqrt(6291) = 79
"001001111",  -- sqrt(6292) = 79
"001001111",  -- sqrt(6293) = 79
"001001111",  -- sqrt(6294) = 79
"001001111",  -- sqrt(6295) = 79
"001001111",  -- sqrt(6296) = 79
"001001111",  -- sqrt(6297) = 79
"001001111",  -- sqrt(6298) = 79
"001001111",  -- sqrt(6299) = 79
"001001111",  -- sqrt(6300) = 79
"001001111",  -- sqrt(6301) = 79
"001001111",  -- sqrt(6302) = 79
"001001111",  -- sqrt(6303) = 79
"001001111",  -- sqrt(6304) = 79
"001001111",  -- sqrt(6305) = 79
"001001111",  -- sqrt(6306) = 79
"001001111",  -- sqrt(6307) = 79
"001001111",  -- sqrt(6308) = 79
"001001111",  -- sqrt(6309) = 79
"001001111",  -- sqrt(6310) = 79
"001001111",  -- sqrt(6311) = 79
"001001111",  -- sqrt(6312) = 79
"001001111",  -- sqrt(6313) = 79
"001001111",  -- sqrt(6314) = 79
"001001111",  -- sqrt(6315) = 79
"001001111",  -- sqrt(6316) = 79
"001001111",  -- sqrt(6317) = 79
"001001111",  -- sqrt(6318) = 79
"001001111",  -- sqrt(6319) = 79
"001001111",  -- sqrt(6320) = 79
"001010000",  -- sqrt(6321) = 80
"001010000",  -- sqrt(6322) = 80
"001010000",  -- sqrt(6323) = 80
"001010000",  -- sqrt(6324) = 80
"001010000",  -- sqrt(6325) = 80
"001010000",  -- sqrt(6326) = 80
"001010000",  -- sqrt(6327) = 80
"001010000",  -- sqrt(6328) = 80
"001010000",  -- sqrt(6329) = 80
"001010000",  -- sqrt(6330) = 80
"001010000",  -- sqrt(6331) = 80
"001010000",  -- sqrt(6332) = 80
"001010000",  -- sqrt(6333) = 80
"001010000",  -- sqrt(6334) = 80
"001010000",  -- sqrt(6335) = 80
"001010000",  -- sqrt(6336) = 80
"001010000",  -- sqrt(6337) = 80
"001010000",  -- sqrt(6338) = 80
"001010000",  -- sqrt(6339) = 80
"001010000",  -- sqrt(6340) = 80
"001010000",  -- sqrt(6341) = 80
"001010000",  -- sqrt(6342) = 80
"001010000",  -- sqrt(6343) = 80
"001010000",  -- sqrt(6344) = 80
"001010000",  -- sqrt(6345) = 80
"001010000",  -- sqrt(6346) = 80
"001010000",  -- sqrt(6347) = 80
"001010000",  -- sqrt(6348) = 80
"001010000",  -- sqrt(6349) = 80
"001010000",  -- sqrt(6350) = 80
"001010000",  -- sqrt(6351) = 80
"001010000",  -- sqrt(6352) = 80
"001010000",  -- sqrt(6353) = 80
"001010000",  -- sqrt(6354) = 80
"001010000",  -- sqrt(6355) = 80
"001010000",  -- sqrt(6356) = 80
"001010000",  -- sqrt(6357) = 80
"001010000",  -- sqrt(6358) = 80
"001010000",  -- sqrt(6359) = 80
"001010000",  -- sqrt(6360) = 80
"001010000",  -- sqrt(6361) = 80
"001010000",  -- sqrt(6362) = 80
"001010000",  -- sqrt(6363) = 80
"001010000",  -- sqrt(6364) = 80
"001010000",  -- sqrt(6365) = 80
"001010000",  -- sqrt(6366) = 80
"001010000",  -- sqrt(6367) = 80
"001010000",  -- sqrt(6368) = 80
"001010000",  -- sqrt(6369) = 80
"001010000",  -- sqrt(6370) = 80
"001010000",  -- sqrt(6371) = 80
"001010000",  -- sqrt(6372) = 80
"001010000",  -- sqrt(6373) = 80
"001010000",  -- sqrt(6374) = 80
"001010000",  -- sqrt(6375) = 80
"001010000",  -- sqrt(6376) = 80
"001010000",  -- sqrt(6377) = 80
"001010000",  -- sqrt(6378) = 80
"001010000",  -- sqrt(6379) = 80
"001010000",  -- sqrt(6380) = 80
"001010000",  -- sqrt(6381) = 80
"001010000",  -- sqrt(6382) = 80
"001010000",  -- sqrt(6383) = 80
"001010000",  -- sqrt(6384) = 80
"001010000",  -- sqrt(6385) = 80
"001010000",  -- sqrt(6386) = 80
"001010000",  -- sqrt(6387) = 80
"001010000",  -- sqrt(6388) = 80
"001010000",  -- sqrt(6389) = 80
"001010000",  -- sqrt(6390) = 80
"001010000",  -- sqrt(6391) = 80
"001010000",  -- sqrt(6392) = 80
"001010000",  -- sqrt(6393) = 80
"001010000",  -- sqrt(6394) = 80
"001010000",  -- sqrt(6395) = 80
"001010000",  -- sqrt(6396) = 80
"001010000",  -- sqrt(6397) = 80
"001010000",  -- sqrt(6398) = 80
"001010000",  -- sqrt(6399) = 80
"001010000",  -- sqrt(6400) = 80
"001010000",  -- sqrt(6401) = 80
"001010000",  -- sqrt(6402) = 80
"001010000",  -- sqrt(6403) = 80
"001010000",  -- sqrt(6404) = 80
"001010000",  -- sqrt(6405) = 80
"001010000",  -- sqrt(6406) = 80
"001010000",  -- sqrt(6407) = 80
"001010000",  -- sqrt(6408) = 80
"001010000",  -- sqrt(6409) = 80
"001010000",  -- sqrt(6410) = 80
"001010000",  -- sqrt(6411) = 80
"001010000",  -- sqrt(6412) = 80
"001010000",  -- sqrt(6413) = 80
"001010000",  -- sqrt(6414) = 80
"001010000",  -- sqrt(6415) = 80
"001010000",  -- sqrt(6416) = 80
"001010000",  -- sqrt(6417) = 80
"001010000",  -- sqrt(6418) = 80
"001010000",  -- sqrt(6419) = 80
"001010000",  -- sqrt(6420) = 80
"001010000",  -- sqrt(6421) = 80
"001010000",  -- sqrt(6422) = 80
"001010000",  -- sqrt(6423) = 80
"001010000",  -- sqrt(6424) = 80
"001010000",  -- sqrt(6425) = 80
"001010000",  -- sqrt(6426) = 80
"001010000",  -- sqrt(6427) = 80
"001010000",  -- sqrt(6428) = 80
"001010000",  -- sqrt(6429) = 80
"001010000",  -- sqrt(6430) = 80
"001010000",  -- sqrt(6431) = 80
"001010000",  -- sqrt(6432) = 80
"001010000",  -- sqrt(6433) = 80
"001010000",  -- sqrt(6434) = 80
"001010000",  -- sqrt(6435) = 80
"001010000",  -- sqrt(6436) = 80
"001010000",  -- sqrt(6437) = 80
"001010000",  -- sqrt(6438) = 80
"001010000",  -- sqrt(6439) = 80
"001010000",  -- sqrt(6440) = 80
"001010000",  -- sqrt(6441) = 80
"001010000",  -- sqrt(6442) = 80
"001010000",  -- sqrt(6443) = 80
"001010000",  -- sqrt(6444) = 80
"001010000",  -- sqrt(6445) = 80
"001010000",  -- sqrt(6446) = 80
"001010000",  -- sqrt(6447) = 80
"001010000",  -- sqrt(6448) = 80
"001010000",  -- sqrt(6449) = 80
"001010000",  -- sqrt(6450) = 80
"001010000",  -- sqrt(6451) = 80
"001010000",  -- sqrt(6452) = 80
"001010000",  -- sqrt(6453) = 80
"001010000",  -- sqrt(6454) = 80
"001010000",  -- sqrt(6455) = 80
"001010000",  -- sqrt(6456) = 80
"001010000",  -- sqrt(6457) = 80
"001010000",  -- sqrt(6458) = 80
"001010000",  -- sqrt(6459) = 80
"001010000",  -- sqrt(6460) = 80
"001010000",  -- sqrt(6461) = 80
"001010000",  -- sqrt(6462) = 80
"001010000",  -- sqrt(6463) = 80
"001010000",  -- sqrt(6464) = 80
"001010000",  -- sqrt(6465) = 80
"001010000",  -- sqrt(6466) = 80
"001010000",  -- sqrt(6467) = 80
"001010000",  -- sqrt(6468) = 80
"001010000",  -- sqrt(6469) = 80
"001010000",  -- sqrt(6470) = 80
"001010000",  -- sqrt(6471) = 80
"001010000",  -- sqrt(6472) = 80
"001010000",  -- sqrt(6473) = 80
"001010000",  -- sqrt(6474) = 80
"001010000",  -- sqrt(6475) = 80
"001010000",  -- sqrt(6476) = 80
"001010000",  -- sqrt(6477) = 80
"001010000",  -- sqrt(6478) = 80
"001010000",  -- sqrt(6479) = 80
"001010000",  -- sqrt(6480) = 80
"001010001",  -- sqrt(6481) = 81
"001010001",  -- sqrt(6482) = 81
"001010001",  -- sqrt(6483) = 81
"001010001",  -- sqrt(6484) = 81
"001010001",  -- sqrt(6485) = 81
"001010001",  -- sqrt(6486) = 81
"001010001",  -- sqrt(6487) = 81
"001010001",  -- sqrt(6488) = 81
"001010001",  -- sqrt(6489) = 81
"001010001",  -- sqrt(6490) = 81
"001010001",  -- sqrt(6491) = 81
"001010001",  -- sqrt(6492) = 81
"001010001",  -- sqrt(6493) = 81
"001010001",  -- sqrt(6494) = 81
"001010001",  -- sqrt(6495) = 81
"001010001",  -- sqrt(6496) = 81
"001010001",  -- sqrt(6497) = 81
"001010001",  -- sqrt(6498) = 81
"001010001",  -- sqrt(6499) = 81
"001010001",  -- sqrt(6500) = 81
"001010001",  -- sqrt(6501) = 81
"001010001",  -- sqrt(6502) = 81
"001010001",  -- sqrt(6503) = 81
"001010001",  -- sqrt(6504) = 81
"001010001",  -- sqrt(6505) = 81
"001010001",  -- sqrt(6506) = 81
"001010001",  -- sqrt(6507) = 81
"001010001",  -- sqrt(6508) = 81
"001010001",  -- sqrt(6509) = 81
"001010001",  -- sqrt(6510) = 81
"001010001",  -- sqrt(6511) = 81
"001010001",  -- sqrt(6512) = 81
"001010001",  -- sqrt(6513) = 81
"001010001",  -- sqrt(6514) = 81
"001010001",  -- sqrt(6515) = 81
"001010001",  -- sqrt(6516) = 81
"001010001",  -- sqrt(6517) = 81
"001010001",  -- sqrt(6518) = 81
"001010001",  -- sqrt(6519) = 81
"001010001",  -- sqrt(6520) = 81
"001010001",  -- sqrt(6521) = 81
"001010001",  -- sqrt(6522) = 81
"001010001",  -- sqrt(6523) = 81
"001010001",  -- sqrt(6524) = 81
"001010001",  -- sqrt(6525) = 81
"001010001",  -- sqrt(6526) = 81
"001010001",  -- sqrt(6527) = 81
"001010001",  -- sqrt(6528) = 81
"001010001",  -- sqrt(6529) = 81
"001010001",  -- sqrt(6530) = 81
"001010001",  -- sqrt(6531) = 81
"001010001",  -- sqrt(6532) = 81
"001010001",  -- sqrt(6533) = 81
"001010001",  -- sqrt(6534) = 81
"001010001",  -- sqrt(6535) = 81
"001010001",  -- sqrt(6536) = 81
"001010001",  -- sqrt(6537) = 81
"001010001",  -- sqrt(6538) = 81
"001010001",  -- sqrt(6539) = 81
"001010001",  -- sqrt(6540) = 81
"001010001",  -- sqrt(6541) = 81
"001010001",  -- sqrt(6542) = 81
"001010001",  -- sqrt(6543) = 81
"001010001",  -- sqrt(6544) = 81
"001010001",  -- sqrt(6545) = 81
"001010001",  -- sqrt(6546) = 81
"001010001",  -- sqrt(6547) = 81
"001010001",  -- sqrt(6548) = 81
"001010001",  -- sqrt(6549) = 81
"001010001",  -- sqrt(6550) = 81
"001010001",  -- sqrt(6551) = 81
"001010001",  -- sqrt(6552) = 81
"001010001",  -- sqrt(6553) = 81
"001010001",  -- sqrt(6554) = 81
"001010001",  -- sqrt(6555) = 81
"001010001",  -- sqrt(6556) = 81
"001010001",  -- sqrt(6557) = 81
"001010001",  -- sqrt(6558) = 81
"001010001",  -- sqrt(6559) = 81
"001010001",  -- sqrt(6560) = 81
"001010001",  -- sqrt(6561) = 81
"001010001",  -- sqrt(6562) = 81
"001010001",  -- sqrt(6563) = 81
"001010001",  -- sqrt(6564) = 81
"001010001",  -- sqrt(6565) = 81
"001010001",  -- sqrt(6566) = 81
"001010001",  -- sqrt(6567) = 81
"001010001",  -- sqrt(6568) = 81
"001010001",  -- sqrt(6569) = 81
"001010001",  -- sqrt(6570) = 81
"001010001",  -- sqrt(6571) = 81
"001010001",  -- sqrt(6572) = 81
"001010001",  -- sqrt(6573) = 81
"001010001",  -- sqrt(6574) = 81
"001010001",  -- sqrt(6575) = 81
"001010001",  -- sqrt(6576) = 81
"001010001",  -- sqrt(6577) = 81
"001010001",  -- sqrt(6578) = 81
"001010001",  -- sqrt(6579) = 81
"001010001",  -- sqrt(6580) = 81
"001010001",  -- sqrt(6581) = 81
"001010001",  -- sqrt(6582) = 81
"001010001",  -- sqrt(6583) = 81
"001010001",  -- sqrt(6584) = 81
"001010001",  -- sqrt(6585) = 81
"001010001",  -- sqrt(6586) = 81
"001010001",  -- sqrt(6587) = 81
"001010001",  -- sqrt(6588) = 81
"001010001",  -- sqrt(6589) = 81
"001010001",  -- sqrt(6590) = 81
"001010001",  -- sqrt(6591) = 81
"001010001",  -- sqrt(6592) = 81
"001010001",  -- sqrt(6593) = 81
"001010001",  -- sqrt(6594) = 81
"001010001",  -- sqrt(6595) = 81
"001010001",  -- sqrt(6596) = 81
"001010001",  -- sqrt(6597) = 81
"001010001",  -- sqrt(6598) = 81
"001010001",  -- sqrt(6599) = 81
"001010001",  -- sqrt(6600) = 81
"001010001",  -- sqrt(6601) = 81
"001010001",  -- sqrt(6602) = 81
"001010001",  -- sqrt(6603) = 81
"001010001",  -- sqrt(6604) = 81
"001010001",  -- sqrt(6605) = 81
"001010001",  -- sqrt(6606) = 81
"001010001",  -- sqrt(6607) = 81
"001010001",  -- sqrt(6608) = 81
"001010001",  -- sqrt(6609) = 81
"001010001",  -- sqrt(6610) = 81
"001010001",  -- sqrt(6611) = 81
"001010001",  -- sqrt(6612) = 81
"001010001",  -- sqrt(6613) = 81
"001010001",  -- sqrt(6614) = 81
"001010001",  -- sqrt(6615) = 81
"001010001",  -- sqrt(6616) = 81
"001010001",  -- sqrt(6617) = 81
"001010001",  -- sqrt(6618) = 81
"001010001",  -- sqrt(6619) = 81
"001010001",  -- sqrt(6620) = 81
"001010001",  -- sqrt(6621) = 81
"001010001",  -- sqrt(6622) = 81
"001010001",  -- sqrt(6623) = 81
"001010001",  -- sqrt(6624) = 81
"001010001",  -- sqrt(6625) = 81
"001010001",  -- sqrt(6626) = 81
"001010001",  -- sqrt(6627) = 81
"001010001",  -- sqrt(6628) = 81
"001010001",  -- sqrt(6629) = 81
"001010001",  -- sqrt(6630) = 81
"001010001",  -- sqrt(6631) = 81
"001010001",  -- sqrt(6632) = 81
"001010001",  -- sqrt(6633) = 81
"001010001",  -- sqrt(6634) = 81
"001010001",  -- sqrt(6635) = 81
"001010001",  -- sqrt(6636) = 81
"001010001",  -- sqrt(6637) = 81
"001010001",  -- sqrt(6638) = 81
"001010001",  -- sqrt(6639) = 81
"001010001",  -- sqrt(6640) = 81
"001010001",  -- sqrt(6641) = 81
"001010001",  -- sqrt(6642) = 81
"001010010",  -- sqrt(6643) = 82
"001010010",  -- sqrt(6644) = 82
"001010010",  -- sqrt(6645) = 82
"001010010",  -- sqrt(6646) = 82
"001010010",  -- sqrt(6647) = 82
"001010010",  -- sqrt(6648) = 82
"001010010",  -- sqrt(6649) = 82
"001010010",  -- sqrt(6650) = 82
"001010010",  -- sqrt(6651) = 82
"001010010",  -- sqrt(6652) = 82
"001010010",  -- sqrt(6653) = 82
"001010010",  -- sqrt(6654) = 82
"001010010",  -- sqrt(6655) = 82
"001010010",  -- sqrt(6656) = 82
"001010010",  -- sqrt(6657) = 82
"001010010",  -- sqrt(6658) = 82
"001010010",  -- sqrt(6659) = 82
"001010010",  -- sqrt(6660) = 82
"001010010",  -- sqrt(6661) = 82
"001010010",  -- sqrt(6662) = 82
"001010010",  -- sqrt(6663) = 82
"001010010",  -- sqrt(6664) = 82
"001010010",  -- sqrt(6665) = 82
"001010010",  -- sqrt(6666) = 82
"001010010",  -- sqrt(6667) = 82
"001010010",  -- sqrt(6668) = 82
"001010010",  -- sqrt(6669) = 82
"001010010",  -- sqrt(6670) = 82
"001010010",  -- sqrt(6671) = 82
"001010010",  -- sqrt(6672) = 82
"001010010",  -- sqrt(6673) = 82
"001010010",  -- sqrt(6674) = 82
"001010010",  -- sqrt(6675) = 82
"001010010",  -- sqrt(6676) = 82
"001010010",  -- sqrt(6677) = 82
"001010010",  -- sqrt(6678) = 82
"001010010",  -- sqrt(6679) = 82
"001010010",  -- sqrt(6680) = 82
"001010010",  -- sqrt(6681) = 82
"001010010",  -- sqrt(6682) = 82
"001010010",  -- sqrt(6683) = 82
"001010010",  -- sqrt(6684) = 82
"001010010",  -- sqrt(6685) = 82
"001010010",  -- sqrt(6686) = 82
"001010010",  -- sqrt(6687) = 82
"001010010",  -- sqrt(6688) = 82
"001010010",  -- sqrt(6689) = 82
"001010010",  -- sqrt(6690) = 82
"001010010",  -- sqrt(6691) = 82
"001010010",  -- sqrt(6692) = 82
"001010010",  -- sqrt(6693) = 82
"001010010",  -- sqrt(6694) = 82
"001010010",  -- sqrt(6695) = 82
"001010010",  -- sqrt(6696) = 82
"001010010",  -- sqrt(6697) = 82
"001010010",  -- sqrt(6698) = 82
"001010010",  -- sqrt(6699) = 82
"001010010",  -- sqrt(6700) = 82
"001010010",  -- sqrt(6701) = 82
"001010010",  -- sqrt(6702) = 82
"001010010",  -- sqrt(6703) = 82
"001010010",  -- sqrt(6704) = 82
"001010010",  -- sqrt(6705) = 82
"001010010",  -- sqrt(6706) = 82
"001010010",  -- sqrt(6707) = 82
"001010010",  -- sqrt(6708) = 82
"001010010",  -- sqrt(6709) = 82
"001010010",  -- sqrt(6710) = 82
"001010010",  -- sqrt(6711) = 82
"001010010",  -- sqrt(6712) = 82
"001010010",  -- sqrt(6713) = 82
"001010010",  -- sqrt(6714) = 82
"001010010",  -- sqrt(6715) = 82
"001010010",  -- sqrt(6716) = 82
"001010010",  -- sqrt(6717) = 82
"001010010",  -- sqrt(6718) = 82
"001010010",  -- sqrt(6719) = 82
"001010010",  -- sqrt(6720) = 82
"001010010",  -- sqrt(6721) = 82
"001010010",  -- sqrt(6722) = 82
"001010010",  -- sqrt(6723) = 82
"001010010",  -- sqrt(6724) = 82
"001010010",  -- sqrt(6725) = 82
"001010010",  -- sqrt(6726) = 82
"001010010",  -- sqrt(6727) = 82
"001010010",  -- sqrt(6728) = 82
"001010010",  -- sqrt(6729) = 82
"001010010",  -- sqrt(6730) = 82
"001010010",  -- sqrt(6731) = 82
"001010010",  -- sqrt(6732) = 82
"001010010",  -- sqrt(6733) = 82
"001010010",  -- sqrt(6734) = 82
"001010010",  -- sqrt(6735) = 82
"001010010",  -- sqrt(6736) = 82
"001010010",  -- sqrt(6737) = 82
"001010010",  -- sqrt(6738) = 82
"001010010",  -- sqrt(6739) = 82
"001010010",  -- sqrt(6740) = 82
"001010010",  -- sqrt(6741) = 82
"001010010",  -- sqrt(6742) = 82
"001010010",  -- sqrt(6743) = 82
"001010010",  -- sqrt(6744) = 82
"001010010",  -- sqrt(6745) = 82
"001010010",  -- sqrt(6746) = 82
"001010010",  -- sqrt(6747) = 82
"001010010",  -- sqrt(6748) = 82
"001010010",  -- sqrt(6749) = 82
"001010010",  -- sqrt(6750) = 82
"001010010",  -- sqrt(6751) = 82
"001010010",  -- sqrt(6752) = 82
"001010010",  -- sqrt(6753) = 82
"001010010",  -- sqrt(6754) = 82
"001010010",  -- sqrt(6755) = 82
"001010010",  -- sqrt(6756) = 82
"001010010",  -- sqrt(6757) = 82
"001010010",  -- sqrt(6758) = 82
"001010010",  -- sqrt(6759) = 82
"001010010",  -- sqrt(6760) = 82
"001010010",  -- sqrt(6761) = 82
"001010010",  -- sqrt(6762) = 82
"001010010",  -- sqrt(6763) = 82
"001010010",  -- sqrt(6764) = 82
"001010010",  -- sqrt(6765) = 82
"001010010",  -- sqrt(6766) = 82
"001010010",  -- sqrt(6767) = 82
"001010010",  -- sqrt(6768) = 82
"001010010",  -- sqrt(6769) = 82
"001010010",  -- sqrt(6770) = 82
"001010010",  -- sqrt(6771) = 82
"001010010",  -- sqrt(6772) = 82
"001010010",  -- sqrt(6773) = 82
"001010010",  -- sqrt(6774) = 82
"001010010",  -- sqrt(6775) = 82
"001010010",  -- sqrt(6776) = 82
"001010010",  -- sqrt(6777) = 82
"001010010",  -- sqrt(6778) = 82
"001010010",  -- sqrt(6779) = 82
"001010010",  -- sqrt(6780) = 82
"001010010",  -- sqrt(6781) = 82
"001010010",  -- sqrt(6782) = 82
"001010010",  -- sqrt(6783) = 82
"001010010",  -- sqrt(6784) = 82
"001010010",  -- sqrt(6785) = 82
"001010010",  -- sqrt(6786) = 82
"001010010",  -- sqrt(6787) = 82
"001010010",  -- sqrt(6788) = 82
"001010010",  -- sqrt(6789) = 82
"001010010",  -- sqrt(6790) = 82
"001010010",  -- sqrt(6791) = 82
"001010010",  -- sqrt(6792) = 82
"001010010",  -- sqrt(6793) = 82
"001010010",  -- sqrt(6794) = 82
"001010010",  -- sqrt(6795) = 82
"001010010",  -- sqrt(6796) = 82
"001010010",  -- sqrt(6797) = 82
"001010010",  -- sqrt(6798) = 82
"001010010",  -- sqrt(6799) = 82
"001010010",  -- sqrt(6800) = 82
"001010010",  -- sqrt(6801) = 82
"001010010",  -- sqrt(6802) = 82
"001010010",  -- sqrt(6803) = 82
"001010010",  -- sqrt(6804) = 82
"001010010",  -- sqrt(6805) = 82
"001010010",  -- sqrt(6806) = 82
"001010011",  -- sqrt(6807) = 83
"001010011",  -- sqrt(6808) = 83
"001010011",  -- sqrt(6809) = 83
"001010011",  -- sqrt(6810) = 83
"001010011",  -- sqrt(6811) = 83
"001010011",  -- sqrt(6812) = 83
"001010011",  -- sqrt(6813) = 83
"001010011",  -- sqrt(6814) = 83
"001010011",  -- sqrt(6815) = 83
"001010011",  -- sqrt(6816) = 83
"001010011",  -- sqrt(6817) = 83
"001010011",  -- sqrt(6818) = 83
"001010011",  -- sqrt(6819) = 83
"001010011",  -- sqrt(6820) = 83
"001010011",  -- sqrt(6821) = 83
"001010011",  -- sqrt(6822) = 83
"001010011",  -- sqrt(6823) = 83
"001010011",  -- sqrt(6824) = 83
"001010011",  -- sqrt(6825) = 83
"001010011",  -- sqrt(6826) = 83
"001010011",  -- sqrt(6827) = 83
"001010011",  -- sqrt(6828) = 83
"001010011",  -- sqrt(6829) = 83
"001010011",  -- sqrt(6830) = 83
"001010011",  -- sqrt(6831) = 83
"001010011",  -- sqrt(6832) = 83
"001010011",  -- sqrt(6833) = 83
"001010011",  -- sqrt(6834) = 83
"001010011",  -- sqrt(6835) = 83
"001010011",  -- sqrt(6836) = 83
"001010011",  -- sqrt(6837) = 83
"001010011",  -- sqrt(6838) = 83
"001010011",  -- sqrt(6839) = 83
"001010011",  -- sqrt(6840) = 83
"001010011",  -- sqrt(6841) = 83
"001010011",  -- sqrt(6842) = 83
"001010011",  -- sqrt(6843) = 83
"001010011",  -- sqrt(6844) = 83
"001010011",  -- sqrt(6845) = 83
"001010011",  -- sqrt(6846) = 83
"001010011",  -- sqrt(6847) = 83
"001010011",  -- sqrt(6848) = 83
"001010011",  -- sqrt(6849) = 83
"001010011",  -- sqrt(6850) = 83
"001010011",  -- sqrt(6851) = 83
"001010011",  -- sqrt(6852) = 83
"001010011",  -- sqrt(6853) = 83
"001010011",  -- sqrt(6854) = 83
"001010011",  -- sqrt(6855) = 83
"001010011",  -- sqrt(6856) = 83
"001010011",  -- sqrt(6857) = 83
"001010011",  -- sqrt(6858) = 83
"001010011",  -- sqrt(6859) = 83
"001010011",  -- sqrt(6860) = 83
"001010011",  -- sqrt(6861) = 83
"001010011",  -- sqrt(6862) = 83
"001010011",  -- sqrt(6863) = 83
"001010011",  -- sqrt(6864) = 83
"001010011",  -- sqrt(6865) = 83
"001010011",  -- sqrt(6866) = 83
"001010011",  -- sqrt(6867) = 83
"001010011",  -- sqrt(6868) = 83
"001010011",  -- sqrt(6869) = 83
"001010011",  -- sqrt(6870) = 83
"001010011",  -- sqrt(6871) = 83
"001010011",  -- sqrt(6872) = 83
"001010011",  -- sqrt(6873) = 83
"001010011",  -- sqrt(6874) = 83
"001010011",  -- sqrt(6875) = 83
"001010011",  -- sqrt(6876) = 83
"001010011",  -- sqrt(6877) = 83
"001010011",  -- sqrt(6878) = 83
"001010011",  -- sqrt(6879) = 83
"001010011",  -- sqrt(6880) = 83
"001010011",  -- sqrt(6881) = 83
"001010011",  -- sqrt(6882) = 83
"001010011",  -- sqrt(6883) = 83
"001010011",  -- sqrt(6884) = 83
"001010011",  -- sqrt(6885) = 83
"001010011",  -- sqrt(6886) = 83
"001010011",  -- sqrt(6887) = 83
"001010011",  -- sqrt(6888) = 83
"001010011",  -- sqrt(6889) = 83
"001010011",  -- sqrt(6890) = 83
"001010011",  -- sqrt(6891) = 83
"001010011",  -- sqrt(6892) = 83
"001010011",  -- sqrt(6893) = 83
"001010011",  -- sqrt(6894) = 83
"001010011",  -- sqrt(6895) = 83
"001010011",  -- sqrt(6896) = 83
"001010011",  -- sqrt(6897) = 83
"001010011",  -- sqrt(6898) = 83
"001010011",  -- sqrt(6899) = 83
"001010011",  -- sqrt(6900) = 83
"001010011",  -- sqrt(6901) = 83
"001010011",  -- sqrt(6902) = 83
"001010011",  -- sqrt(6903) = 83
"001010011",  -- sqrt(6904) = 83
"001010011",  -- sqrt(6905) = 83
"001010011",  -- sqrt(6906) = 83
"001010011",  -- sqrt(6907) = 83
"001010011",  -- sqrt(6908) = 83
"001010011",  -- sqrt(6909) = 83
"001010011",  -- sqrt(6910) = 83
"001010011",  -- sqrt(6911) = 83
"001010011",  -- sqrt(6912) = 83
"001010011",  -- sqrt(6913) = 83
"001010011",  -- sqrt(6914) = 83
"001010011",  -- sqrt(6915) = 83
"001010011",  -- sqrt(6916) = 83
"001010011",  -- sqrt(6917) = 83
"001010011",  -- sqrt(6918) = 83
"001010011",  -- sqrt(6919) = 83
"001010011",  -- sqrt(6920) = 83
"001010011",  -- sqrt(6921) = 83
"001010011",  -- sqrt(6922) = 83
"001010011",  -- sqrt(6923) = 83
"001010011",  -- sqrt(6924) = 83
"001010011",  -- sqrt(6925) = 83
"001010011",  -- sqrt(6926) = 83
"001010011",  -- sqrt(6927) = 83
"001010011",  -- sqrt(6928) = 83
"001010011",  -- sqrt(6929) = 83
"001010011",  -- sqrt(6930) = 83
"001010011",  -- sqrt(6931) = 83
"001010011",  -- sqrt(6932) = 83
"001010011",  -- sqrt(6933) = 83
"001010011",  -- sqrt(6934) = 83
"001010011",  -- sqrt(6935) = 83
"001010011",  -- sqrt(6936) = 83
"001010011",  -- sqrt(6937) = 83
"001010011",  -- sqrt(6938) = 83
"001010011",  -- sqrt(6939) = 83
"001010011",  -- sqrt(6940) = 83
"001010011",  -- sqrt(6941) = 83
"001010011",  -- sqrt(6942) = 83
"001010011",  -- sqrt(6943) = 83
"001010011",  -- sqrt(6944) = 83
"001010011",  -- sqrt(6945) = 83
"001010011",  -- sqrt(6946) = 83
"001010011",  -- sqrt(6947) = 83
"001010011",  -- sqrt(6948) = 83
"001010011",  -- sqrt(6949) = 83
"001010011",  -- sqrt(6950) = 83
"001010011",  -- sqrt(6951) = 83
"001010011",  -- sqrt(6952) = 83
"001010011",  -- sqrt(6953) = 83
"001010011",  -- sqrt(6954) = 83
"001010011",  -- sqrt(6955) = 83
"001010011",  -- sqrt(6956) = 83
"001010011",  -- sqrt(6957) = 83
"001010011",  -- sqrt(6958) = 83
"001010011",  -- sqrt(6959) = 83
"001010011",  -- sqrt(6960) = 83
"001010011",  -- sqrt(6961) = 83
"001010011",  -- sqrt(6962) = 83
"001010011",  -- sqrt(6963) = 83
"001010011",  -- sqrt(6964) = 83
"001010011",  -- sqrt(6965) = 83
"001010011",  -- sqrt(6966) = 83
"001010011",  -- sqrt(6967) = 83
"001010011",  -- sqrt(6968) = 83
"001010011",  -- sqrt(6969) = 83
"001010011",  -- sqrt(6970) = 83
"001010011",  -- sqrt(6971) = 83
"001010011",  -- sqrt(6972) = 83
"001010100",  -- sqrt(6973) = 84
"001010100",  -- sqrt(6974) = 84
"001010100",  -- sqrt(6975) = 84
"001010100",  -- sqrt(6976) = 84
"001010100",  -- sqrt(6977) = 84
"001010100",  -- sqrt(6978) = 84
"001010100",  -- sqrt(6979) = 84
"001010100",  -- sqrt(6980) = 84
"001010100",  -- sqrt(6981) = 84
"001010100",  -- sqrt(6982) = 84
"001010100",  -- sqrt(6983) = 84
"001010100",  -- sqrt(6984) = 84
"001010100",  -- sqrt(6985) = 84
"001010100",  -- sqrt(6986) = 84
"001010100",  -- sqrt(6987) = 84
"001010100",  -- sqrt(6988) = 84
"001010100",  -- sqrt(6989) = 84
"001010100",  -- sqrt(6990) = 84
"001010100",  -- sqrt(6991) = 84
"001010100",  -- sqrt(6992) = 84
"001010100",  -- sqrt(6993) = 84
"001010100",  -- sqrt(6994) = 84
"001010100",  -- sqrt(6995) = 84
"001010100",  -- sqrt(6996) = 84
"001010100",  -- sqrt(6997) = 84
"001010100",  -- sqrt(6998) = 84
"001010100",  -- sqrt(6999) = 84
"001010100",  -- sqrt(7000) = 84
"001010100",  -- sqrt(7001) = 84
"001010100",  -- sqrt(7002) = 84
"001010100",  -- sqrt(7003) = 84
"001010100",  -- sqrt(7004) = 84
"001010100",  -- sqrt(7005) = 84
"001010100",  -- sqrt(7006) = 84
"001010100",  -- sqrt(7007) = 84
"001010100",  -- sqrt(7008) = 84
"001010100",  -- sqrt(7009) = 84
"001010100",  -- sqrt(7010) = 84
"001010100",  -- sqrt(7011) = 84
"001010100",  -- sqrt(7012) = 84
"001010100",  -- sqrt(7013) = 84
"001010100",  -- sqrt(7014) = 84
"001010100",  -- sqrt(7015) = 84
"001010100",  -- sqrt(7016) = 84
"001010100",  -- sqrt(7017) = 84
"001010100",  -- sqrt(7018) = 84
"001010100",  -- sqrt(7019) = 84
"001010100",  -- sqrt(7020) = 84
"001010100",  -- sqrt(7021) = 84
"001010100",  -- sqrt(7022) = 84
"001010100",  -- sqrt(7023) = 84
"001010100",  -- sqrt(7024) = 84
"001010100",  -- sqrt(7025) = 84
"001010100",  -- sqrt(7026) = 84
"001010100",  -- sqrt(7027) = 84
"001010100",  -- sqrt(7028) = 84
"001010100",  -- sqrt(7029) = 84
"001010100",  -- sqrt(7030) = 84
"001010100",  -- sqrt(7031) = 84
"001010100",  -- sqrt(7032) = 84
"001010100",  -- sqrt(7033) = 84
"001010100",  -- sqrt(7034) = 84
"001010100",  -- sqrt(7035) = 84
"001010100",  -- sqrt(7036) = 84
"001010100",  -- sqrt(7037) = 84
"001010100",  -- sqrt(7038) = 84
"001010100",  -- sqrt(7039) = 84
"001010100",  -- sqrt(7040) = 84
"001010100",  -- sqrt(7041) = 84
"001010100",  -- sqrt(7042) = 84
"001010100",  -- sqrt(7043) = 84
"001010100",  -- sqrt(7044) = 84
"001010100",  -- sqrt(7045) = 84
"001010100",  -- sqrt(7046) = 84
"001010100",  -- sqrt(7047) = 84
"001010100",  -- sqrt(7048) = 84
"001010100",  -- sqrt(7049) = 84
"001010100",  -- sqrt(7050) = 84
"001010100",  -- sqrt(7051) = 84
"001010100",  -- sqrt(7052) = 84
"001010100",  -- sqrt(7053) = 84
"001010100",  -- sqrt(7054) = 84
"001010100",  -- sqrt(7055) = 84
"001010100",  -- sqrt(7056) = 84
"001010100",  -- sqrt(7057) = 84
"001010100",  -- sqrt(7058) = 84
"001010100",  -- sqrt(7059) = 84
"001010100",  -- sqrt(7060) = 84
"001010100",  -- sqrt(7061) = 84
"001010100",  -- sqrt(7062) = 84
"001010100",  -- sqrt(7063) = 84
"001010100",  -- sqrt(7064) = 84
"001010100",  -- sqrt(7065) = 84
"001010100",  -- sqrt(7066) = 84
"001010100",  -- sqrt(7067) = 84
"001010100",  -- sqrt(7068) = 84
"001010100",  -- sqrt(7069) = 84
"001010100",  -- sqrt(7070) = 84
"001010100",  -- sqrt(7071) = 84
"001010100",  -- sqrt(7072) = 84
"001010100",  -- sqrt(7073) = 84
"001010100",  -- sqrt(7074) = 84
"001010100",  -- sqrt(7075) = 84
"001010100",  -- sqrt(7076) = 84
"001010100",  -- sqrt(7077) = 84
"001010100",  -- sqrt(7078) = 84
"001010100",  -- sqrt(7079) = 84
"001010100",  -- sqrt(7080) = 84
"001010100",  -- sqrt(7081) = 84
"001010100",  -- sqrt(7082) = 84
"001010100",  -- sqrt(7083) = 84
"001010100",  -- sqrt(7084) = 84
"001010100",  -- sqrt(7085) = 84
"001010100",  -- sqrt(7086) = 84
"001010100",  -- sqrt(7087) = 84
"001010100",  -- sqrt(7088) = 84
"001010100",  -- sqrt(7089) = 84
"001010100",  -- sqrt(7090) = 84
"001010100",  -- sqrt(7091) = 84
"001010100",  -- sqrt(7092) = 84
"001010100",  -- sqrt(7093) = 84
"001010100",  -- sqrt(7094) = 84
"001010100",  -- sqrt(7095) = 84
"001010100",  -- sqrt(7096) = 84
"001010100",  -- sqrt(7097) = 84
"001010100",  -- sqrt(7098) = 84
"001010100",  -- sqrt(7099) = 84
"001010100",  -- sqrt(7100) = 84
"001010100",  -- sqrt(7101) = 84
"001010100",  -- sqrt(7102) = 84
"001010100",  -- sqrt(7103) = 84
"001010100",  -- sqrt(7104) = 84
"001010100",  -- sqrt(7105) = 84
"001010100",  -- sqrt(7106) = 84
"001010100",  -- sqrt(7107) = 84
"001010100",  -- sqrt(7108) = 84
"001010100",  -- sqrt(7109) = 84
"001010100",  -- sqrt(7110) = 84
"001010100",  -- sqrt(7111) = 84
"001010100",  -- sqrt(7112) = 84
"001010100",  -- sqrt(7113) = 84
"001010100",  -- sqrt(7114) = 84
"001010100",  -- sqrt(7115) = 84
"001010100",  -- sqrt(7116) = 84
"001010100",  -- sqrt(7117) = 84
"001010100",  -- sqrt(7118) = 84
"001010100",  -- sqrt(7119) = 84
"001010100",  -- sqrt(7120) = 84
"001010100",  -- sqrt(7121) = 84
"001010100",  -- sqrt(7122) = 84
"001010100",  -- sqrt(7123) = 84
"001010100",  -- sqrt(7124) = 84
"001010100",  -- sqrt(7125) = 84
"001010100",  -- sqrt(7126) = 84
"001010100",  -- sqrt(7127) = 84
"001010100",  -- sqrt(7128) = 84
"001010100",  -- sqrt(7129) = 84
"001010100",  -- sqrt(7130) = 84
"001010100",  -- sqrt(7131) = 84
"001010100",  -- sqrt(7132) = 84
"001010100",  -- sqrt(7133) = 84
"001010100",  -- sqrt(7134) = 84
"001010100",  -- sqrt(7135) = 84
"001010100",  -- sqrt(7136) = 84
"001010100",  -- sqrt(7137) = 84
"001010100",  -- sqrt(7138) = 84
"001010100",  -- sqrt(7139) = 84
"001010100",  -- sqrt(7140) = 84
"001010101",  -- sqrt(7141) = 85
"001010101",  -- sqrt(7142) = 85
"001010101",  -- sqrt(7143) = 85
"001010101",  -- sqrt(7144) = 85
"001010101",  -- sqrt(7145) = 85
"001010101",  -- sqrt(7146) = 85
"001010101",  -- sqrt(7147) = 85
"001010101",  -- sqrt(7148) = 85
"001010101",  -- sqrt(7149) = 85
"001010101",  -- sqrt(7150) = 85
"001010101",  -- sqrt(7151) = 85
"001010101",  -- sqrt(7152) = 85
"001010101",  -- sqrt(7153) = 85
"001010101",  -- sqrt(7154) = 85
"001010101",  -- sqrt(7155) = 85
"001010101",  -- sqrt(7156) = 85
"001010101",  -- sqrt(7157) = 85
"001010101",  -- sqrt(7158) = 85
"001010101",  -- sqrt(7159) = 85
"001010101",  -- sqrt(7160) = 85
"001010101",  -- sqrt(7161) = 85
"001010101",  -- sqrt(7162) = 85
"001010101",  -- sqrt(7163) = 85
"001010101",  -- sqrt(7164) = 85
"001010101",  -- sqrt(7165) = 85
"001010101",  -- sqrt(7166) = 85
"001010101",  -- sqrt(7167) = 85
"001010101",  -- sqrt(7168) = 85
"001010101",  -- sqrt(7169) = 85
"001010101",  -- sqrt(7170) = 85
"001010101",  -- sqrt(7171) = 85
"001010101",  -- sqrt(7172) = 85
"001010101",  -- sqrt(7173) = 85
"001010101",  -- sqrt(7174) = 85
"001010101",  -- sqrt(7175) = 85
"001010101",  -- sqrt(7176) = 85
"001010101",  -- sqrt(7177) = 85
"001010101",  -- sqrt(7178) = 85
"001010101",  -- sqrt(7179) = 85
"001010101",  -- sqrt(7180) = 85
"001010101",  -- sqrt(7181) = 85
"001010101",  -- sqrt(7182) = 85
"001010101",  -- sqrt(7183) = 85
"001010101",  -- sqrt(7184) = 85
"001010101",  -- sqrt(7185) = 85
"001010101",  -- sqrt(7186) = 85
"001010101",  -- sqrt(7187) = 85
"001010101",  -- sqrt(7188) = 85
"001010101",  -- sqrt(7189) = 85
"001010101",  -- sqrt(7190) = 85
"001010101",  -- sqrt(7191) = 85
"001010101",  -- sqrt(7192) = 85
"001010101",  -- sqrt(7193) = 85
"001010101",  -- sqrt(7194) = 85
"001010101",  -- sqrt(7195) = 85
"001010101",  -- sqrt(7196) = 85
"001010101",  -- sqrt(7197) = 85
"001010101",  -- sqrt(7198) = 85
"001010101",  -- sqrt(7199) = 85
"001010101",  -- sqrt(7200) = 85
"001010101",  -- sqrt(7201) = 85
"001010101",  -- sqrt(7202) = 85
"001010101",  -- sqrt(7203) = 85
"001010101",  -- sqrt(7204) = 85
"001010101",  -- sqrt(7205) = 85
"001010101",  -- sqrt(7206) = 85
"001010101",  -- sqrt(7207) = 85
"001010101",  -- sqrt(7208) = 85
"001010101",  -- sqrt(7209) = 85
"001010101",  -- sqrt(7210) = 85
"001010101",  -- sqrt(7211) = 85
"001010101",  -- sqrt(7212) = 85
"001010101",  -- sqrt(7213) = 85
"001010101",  -- sqrt(7214) = 85
"001010101",  -- sqrt(7215) = 85
"001010101",  -- sqrt(7216) = 85
"001010101",  -- sqrt(7217) = 85
"001010101",  -- sqrt(7218) = 85
"001010101",  -- sqrt(7219) = 85
"001010101",  -- sqrt(7220) = 85
"001010101",  -- sqrt(7221) = 85
"001010101",  -- sqrt(7222) = 85
"001010101",  -- sqrt(7223) = 85
"001010101",  -- sqrt(7224) = 85
"001010101",  -- sqrt(7225) = 85
"001010101",  -- sqrt(7226) = 85
"001010101",  -- sqrt(7227) = 85
"001010101",  -- sqrt(7228) = 85
"001010101",  -- sqrt(7229) = 85
"001010101",  -- sqrt(7230) = 85
"001010101",  -- sqrt(7231) = 85
"001010101",  -- sqrt(7232) = 85
"001010101",  -- sqrt(7233) = 85
"001010101",  -- sqrt(7234) = 85
"001010101",  -- sqrt(7235) = 85
"001010101",  -- sqrt(7236) = 85
"001010101",  -- sqrt(7237) = 85
"001010101",  -- sqrt(7238) = 85
"001010101",  -- sqrt(7239) = 85
"001010101",  -- sqrt(7240) = 85
"001010101",  -- sqrt(7241) = 85
"001010101",  -- sqrt(7242) = 85
"001010101",  -- sqrt(7243) = 85
"001010101",  -- sqrt(7244) = 85
"001010101",  -- sqrt(7245) = 85
"001010101",  -- sqrt(7246) = 85
"001010101",  -- sqrt(7247) = 85
"001010101",  -- sqrt(7248) = 85
"001010101",  -- sqrt(7249) = 85
"001010101",  -- sqrt(7250) = 85
"001010101",  -- sqrt(7251) = 85
"001010101",  -- sqrt(7252) = 85
"001010101",  -- sqrt(7253) = 85
"001010101",  -- sqrt(7254) = 85
"001010101",  -- sqrt(7255) = 85
"001010101",  -- sqrt(7256) = 85
"001010101",  -- sqrt(7257) = 85
"001010101",  -- sqrt(7258) = 85
"001010101",  -- sqrt(7259) = 85
"001010101",  -- sqrt(7260) = 85
"001010101",  -- sqrt(7261) = 85
"001010101",  -- sqrt(7262) = 85
"001010101",  -- sqrt(7263) = 85
"001010101",  -- sqrt(7264) = 85
"001010101",  -- sqrt(7265) = 85
"001010101",  -- sqrt(7266) = 85
"001010101",  -- sqrt(7267) = 85
"001010101",  -- sqrt(7268) = 85
"001010101",  -- sqrt(7269) = 85
"001010101",  -- sqrt(7270) = 85
"001010101",  -- sqrt(7271) = 85
"001010101",  -- sqrt(7272) = 85
"001010101",  -- sqrt(7273) = 85
"001010101",  -- sqrt(7274) = 85
"001010101",  -- sqrt(7275) = 85
"001010101",  -- sqrt(7276) = 85
"001010101",  -- sqrt(7277) = 85
"001010101",  -- sqrt(7278) = 85
"001010101",  -- sqrt(7279) = 85
"001010101",  -- sqrt(7280) = 85
"001010101",  -- sqrt(7281) = 85
"001010101",  -- sqrt(7282) = 85
"001010101",  -- sqrt(7283) = 85
"001010101",  -- sqrt(7284) = 85
"001010101",  -- sqrt(7285) = 85
"001010101",  -- sqrt(7286) = 85
"001010101",  -- sqrt(7287) = 85
"001010101",  -- sqrt(7288) = 85
"001010101",  -- sqrt(7289) = 85
"001010101",  -- sqrt(7290) = 85
"001010101",  -- sqrt(7291) = 85
"001010101",  -- sqrt(7292) = 85
"001010101",  -- sqrt(7293) = 85
"001010101",  -- sqrt(7294) = 85
"001010101",  -- sqrt(7295) = 85
"001010101",  -- sqrt(7296) = 85
"001010101",  -- sqrt(7297) = 85
"001010101",  -- sqrt(7298) = 85
"001010101",  -- sqrt(7299) = 85
"001010101",  -- sqrt(7300) = 85
"001010101",  -- sqrt(7301) = 85
"001010101",  -- sqrt(7302) = 85
"001010101",  -- sqrt(7303) = 85
"001010101",  -- sqrt(7304) = 85
"001010101",  -- sqrt(7305) = 85
"001010101",  -- sqrt(7306) = 85
"001010101",  -- sqrt(7307) = 85
"001010101",  -- sqrt(7308) = 85
"001010101",  -- sqrt(7309) = 85
"001010101",  -- sqrt(7310) = 85
"001010110",  -- sqrt(7311) = 86
"001010110",  -- sqrt(7312) = 86
"001010110",  -- sqrt(7313) = 86
"001010110",  -- sqrt(7314) = 86
"001010110",  -- sqrt(7315) = 86
"001010110",  -- sqrt(7316) = 86
"001010110",  -- sqrt(7317) = 86
"001010110",  -- sqrt(7318) = 86
"001010110",  -- sqrt(7319) = 86
"001010110",  -- sqrt(7320) = 86
"001010110",  -- sqrt(7321) = 86
"001010110",  -- sqrt(7322) = 86
"001010110",  -- sqrt(7323) = 86
"001010110",  -- sqrt(7324) = 86
"001010110",  -- sqrt(7325) = 86
"001010110",  -- sqrt(7326) = 86
"001010110",  -- sqrt(7327) = 86
"001010110",  -- sqrt(7328) = 86
"001010110",  -- sqrt(7329) = 86
"001010110",  -- sqrt(7330) = 86
"001010110",  -- sqrt(7331) = 86
"001010110",  -- sqrt(7332) = 86
"001010110",  -- sqrt(7333) = 86
"001010110",  -- sqrt(7334) = 86
"001010110",  -- sqrt(7335) = 86
"001010110",  -- sqrt(7336) = 86
"001010110",  -- sqrt(7337) = 86
"001010110",  -- sqrt(7338) = 86
"001010110",  -- sqrt(7339) = 86
"001010110",  -- sqrt(7340) = 86
"001010110",  -- sqrt(7341) = 86
"001010110",  -- sqrt(7342) = 86
"001010110",  -- sqrt(7343) = 86
"001010110",  -- sqrt(7344) = 86
"001010110",  -- sqrt(7345) = 86
"001010110",  -- sqrt(7346) = 86
"001010110",  -- sqrt(7347) = 86
"001010110",  -- sqrt(7348) = 86
"001010110",  -- sqrt(7349) = 86
"001010110",  -- sqrt(7350) = 86
"001010110",  -- sqrt(7351) = 86
"001010110",  -- sqrt(7352) = 86
"001010110",  -- sqrt(7353) = 86
"001010110",  -- sqrt(7354) = 86
"001010110",  -- sqrt(7355) = 86
"001010110",  -- sqrt(7356) = 86
"001010110",  -- sqrt(7357) = 86
"001010110",  -- sqrt(7358) = 86
"001010110",  -- sqrt(7359) = 86
"001010110",  -- sqrt(7360) = 86
"001010110",  -- sqrt(7361) = 86
"001010110",  -- sqrt(7362) = 86
"001010110",  -- sqrt(7363) = 86
"001010110",  -- sqrt(7364) = 86
"001010110",  -- sqrt(7365) = 86
"001010110",  -- sqrt(7366) = 86
"001010110",  -- sqrt(7367) = 86
"001010110",  -- sqrt(7368) = 86
"001010110",  -- sqrt(7369) = 86
"001010110",  -- sqrt(7370) = 86
"001010110",  -- sqrt(7371) = 86
"001010110",  -- sqrt(7372) = 86
"001010110",  -- sqrt(7373) = 86
"001010110",  -- sqrt(7374) = 86
"001010110",  -- sqrt(7375) = 86
"001010110",  -- sqrt(7376) = 86
"001010110",  -- sqrt(7377) = 86
"001010110",  -- sqrt(7378) = 86
"001010110",  -- sqrt(7379) = 86
"001010110",  -- sqrt(7380) = 86
"001010110",  -- sqrt(7381) = 86
"001010110",  -- sqrt(7382) = 86
"001010110",  -- sqrt(7383) = 86
"001010110",  -- sqrt(7384) = 86
"001010110",  -- sqrt(7385) = 86
"001010110",  -- sqrt(7386) = 86
"001010110",  -- sqrt(7387) = 86
"001010110",  -- sqrt(7388) = 86
"001010110",  -- sqrt(7389) = 86
"001010110",  -- sqrt(7390) = 86
"001010110",  -- sqrt(7391) = 86
"001010110",  -- sqrt(7392) = 86
"001010110",  -- sqrt(7393) = 86
"001010110",  -- sqrt(7394) = 86
"001010110",  -- sqrt(7395) = 86
"001010110",  -- sqrt(7396) = 86
"001010110",  -- sqrt(7397) = 86
"001010110",  -- sqrt(7398) = 86
"001010110",  -- sqrt(7399) = 86
"001010110",  -- sqrt(7400) = 86
"001010110",  -- sqrt(7401) = 86
"001010110",  -- sqrt(7402) = 86
"001010110",  -- sqrt(7403) = 86
"001010110",  -- sqrt(7404) = 86
"001010110",  -- sqrt(7405) = 86
"001010110",  -- sqrt(7406) = 86
"001010110",  -- sqrt(7407) = 86
"001010110",  -- sqrt(7408) = 86
"001010110",  -- sqrt(7409) = 86
"001010110",  -- sqrt(7410) = 86
"001010110",  -- sqrt(7411) = 86
"001010110",  -- sqrt(7412) = 86
"001010110",  -- sqrt(7413) = 86
"001010110",  -- sqrt(7414) = 86
"001010110",  -- sqrt(7415) = 86
"001010110",  -- sqrt(7416) = 86
"001010110",  -- sqrt(7417) = 86
"001010110",  -- sqrt(7418) = 86
"001010110",  -- sqrt(7419) = 86
"001010110",  -- sqrt(7420) = 86
"001010110",  -- sqrt(7421) = 86
"001010110",  -- sqrt(7422) = 86
"001010110",  -- sqrt(7423) = 86
"001010110",  -- sqrt(7424) = 86
"001010110",  -- sqrt(7425) = 86
"001010110",  -- sqrt(7426) = 86
"001010110",  -- sqrt(7427) = 86
"001010110",  -- sqrt(7428) = 86
"001010110",  -- sqrt(7429) = 86
"001010110",  -- sqrt(7430) = 86
"001010110",  -- sqrt(7431) = 86
"001010110",  -- sqrt(7432) = 86
"001010110",  -- sqrt(7433) = 86
"001010110",  -- sqrt(7434) = 86
"001010110",  -- sqrt(7435) = 86
"001010110",  -- sqrt(7436) = 86
"001010110",  -- sqrt(7437) = 86
"001010110",  -- sqrt(7438) = 86
"001010110",  -- sqrt(7439) = 86
"001010110",  -- sqrt(7440) = 86
"001010110",  -- sqrt(7441) = 86
"001010110",  -- sqrt(7442) = 86
"001010110",  -- sqrt(7443) = 86
"001010110",  -- sqrt(7444) = 86
"001010110",  -- sqrt(7445) = 86
"001010110",  -- sqrt(7446) = 86
"001010110",  -- sqrt(7447) = 86
"001010110",  -- sqrt(7448) = 86
"001010110",  -- sqrt(7449) = 86
"001010110",  -- sqrt(7450) = 86
"001010110",  -- sqrt(7451) = 86
"001010110",  -- sqrt(7452) = 86
"001010110",  -- sqrt(7453) = 86
"001010110",  -- sqrt(7454) = 86
"001010110",  -- sqrt(7455) = 86
"001010110",  -- sqrt(7456) = 86
"001010110",  -- sqrt(7457) = 86
"001010110",  -- sqrt(7458) = 86
"001010110",  -- sqrt(7459) = 86
"001010110",  -- sqrt(7460) = 86
"001010110",  -- sqrt(7461) = 86
"001010110",  -- sqrt(7462) = 86
"001010110",  -- sqrt(7463) = 86
"001010110",  -- sqrt(7464) = 86
"001010110",  -- sqrt(7465) = 86
"001010110",  -- sqrt(7466) = 86
"001010110",  -- sqrt(7467) = 86
"001010110",  -- sqrt(7468) = 86
"001010110",  -- sqrt(7469) = 86
"001010110",  -- sqrt(7470) = 86
"001010110",  -- sqrt(7471) = 86
"001010110",  -- sqrt(7472) = 86
"001010110",  -- sqrt(7473) = 86
"001010110",  -- sqrt(7474) = 86
"001010110",  -- sqrt(7475) = 86
"001010110",  -- sqrt(7476) = 86
"001010110",  -- sqrt(7477) = 86
"001010110",  -- sqrt(7478) = 86
"001010110",  -- sqrt(7479) = 86
"001010110",  -- sqrt(7480) = 86
"001010110",  -- sqrt(7481) = 86
"001010110",  -- sqrt(7482) = 86
"001010111",  -- sqrt(7483) = 87
"001010111",  -- sqrt(7484) = 87
"001010111",  -- sqrt(7485) = 87
"001010111",  -- sqrt(7486) = 87
"001010111",  -- sqrt(7487) = 87
"001010111",  -- sqrt(7488) = 87
"001010111",  -- sqrt(7489) = 87
"001010111",  -- sqrt(7490) = 87
"001010111",  -- sqrt(7491) = 87
"001010111",  -- sqrt(7492) = 87
"001010111",  -- sqrt(7493) = 87
"001010111",  -- sqrt(7494) = 87
"001010111",  -- sqrt(7495) = 87
"001010111",  -- sqrt(7496) = 87
"001010111",  -- sqrt(7497) = 87
"001010111",  -- sqrt(7498) = 87
"001010111",  -- sqrt(7499) = 87
"001010111",  -- sqrt(7500) = 87
"001010111",  -- sqrt(7501) = 87
"001010111",  -- sqrt(7502) = 87
"001010111",  -- sqrt(7503) = 87
"001010111",  -- sqrt(7504) = 87
"001010111",  -- sqrt(7505) = 87
"001010111",  -- sqrt(7506) = 87
"001010111",  -- sqrt(7507) = 87
"001010111",  -- sqrt(7508) = 87
"001010111",  -- sqrt(7509) = 87
"001010111",  -- sqrt(7510) = 87
"001010111",  -- sqrt(7511) = 87
"001010111",  -- sqrt(7512) = 87
"001010111",  -- sqrt(7513) = 87
"001010111",  -- sqrt(7514) = 87
"001010111",  -- sqrt(7515) = 87
"001010111",  -- sqrt(7516) = 87
"001010111",  -- sqrt(7517) = 87
"001010111",  -- sqrt(7518) = 87
"001010111",  -- sqrt(7519) = 87
"001010111",  -- sqrt(7520) = 87
"001010111",  -- sqrt(7521) = 87
"001010111",  -- sqrt(7522) = 87
"001010111",  -- sqrt(7523) = 87
"001010111",  -- sqrt(7524) = 87
"001010111",  -- sqrt(7525) = 87
"001010111",  -- sqrt(7526) = 87
"001010111",  -- sqrt(7527) = 87
"001010111",  -- sqrt(7528) = 87
"001010111",  -- sqrt(7529) = 87
"001010111",  -- sqrt(7530) = 87
"001010111",  -- sqrt(7531) = 87
"001010111",  -- sqrt(7532) = 87
"001010111",  -- sqrt(7533) = 87
"001010111",  -- sqrt(7534) = 87
"001010111",  -- sqrt(7535) = 87
"001010111",  -- sqrt(7536) = 87
"001010111",  -- sqrt(7537) = 87
"001010111",  -- sqrt(7538) = 87
"001010111",  -- sqrt(7539) = 87
"001010111",  -- sqrt(7540) = 87
"001010111",  -- sqrt(7541) = 87
"001010111",  -- sqrt(7542) = 87
"001010111",  -- sqrt(7543) = 87
"001010111",  -- sqrt(7544) = 87
"001010111",  -- sqrt(7545) = 87
"001010111",  -- sqrt(7546) = 87
"001010111",  -- sqrt(7547) = 87
"001010111",  -- sqrt(7548) = 87
"001010111",  -- sqrt(7549) = 87
"001010111",  -- sqrt(7550) = 87
"001010111",  -- sqrt(7551) = 87
"001010111",  -- sqrt(7552) = 87
"001010111",  -- sqrt(7553) = 87
"001010111",  -- sqrt(7554) = 87
"001010111",  -- sqrt(7555) = 87
"001010111",  -- sqrt(7556) = 87
"001010111",  -- sqrt(7557) = 87
"001010111",  -- sqrt(7558) = 87
"001010111",  -- sqrt(7559) = 87
"001010111",  -- sqrt(7560) = 87
"001010111",  -- sqrt(7561) = 87
"001010111",  -- sqrt(7562) = 87
"001010111",  -- sqrt(7563) = 87
"001010111",  -- sqrt(7564) = 87
"001010111",  -- sqrt(7565) = 87
"001010111",  -- sqrt(7566) = 87
"001010111",  -- sqrt(7567) = 87
"001010111",  -- sqrt(7568) = 87
"001010111",  -- sqrt(7569) = 87
"001010111",  -- sqrt(7570) = 87
"001010111",  -- sqrt(7571) = 87
"001010111",  -- sqrt(7572) = 87
"001010111",  -- sqrt(7573) = 87
"001010111",  -- sqrt(7574) = 87
"001010111",  -- sqrt(7575) = 87
"001010111",  -- sqrt(7576) = 87
"001010111",  -- sqrt(7577) = 87
"001010111",  -- sqrt(7578) = 87
"001010111",  -- sqrt(7579) = 87
"001010111",  -- sqrt(7580) = 87
"001010111",  -- sqrt(7581) = 87
"001010111",  -- sqrt(7582) = 87
"001010111",  -- sqrt(7583) = 87
"001010111",  -- sqrt(7584) = 87
"001010111",  -- sqrt(7585) = 87
"001010111",  -- sqrt(7586) = 87
"001010111",  -- sqrt(7587) = 87
"001010111",  -- sqrt(7588) = 87
"001010111",  -- sqrt(7589) = 87
"001010111",  -- sqrt(7590) = 87
"001010111",  -- sqrt(7591) = 87
"001010111",  -- sqrt(7592) = 87
"001010111",  -- sqrt(7593) = 87
"001010111",  -- sqrt(7594) = 87
"001010111",  -- sqrt(7595) = 87
"001010111",  -- sqrt(7596) = 87
"001010111",  -- sqrt(7597) = 87
"001010111",  -- sqrt(7598) = 87
"001010111",  -- sqrt(7599) = 87
"001010111",  -- sqrt(7600) = 87
"001010111",  -- sqrt(7601) = 87
"001010111",  -- sqrt(7602) = 87
"001010111",  -- sqrt(7603) = 87
"001010111",  -- sqrt(7604) = 87
"001010111",  -- sqrt(7605) = 87
"001010111",  -- sqrt(7606) = 87
"001010111",  -- sqrt(7607) = 87
"001010111",  -- sqrt(7608) = 87
"001010111",  -- sqrt(7609) = 87
"001010111",  -- sqrt(7610) = 87
"001010111",  -- sqrt(7611) = 87
"001010111",  -- sqrt(7612) = 87
"001010111",  -- sqrt(7613) = 87
"001010111",  -- sqrt(7614) = 87
"001010111",  -- sqrt(7615) = 87
"001010111",  -- sqrt(7616) = 87
"001010111",  -- sqrt(7617) = 87
"001010111",  -- sqrt(7618) = 87
"001010111",  -- sqrt(7619) = 87
"001010111",  -- sqrt(7620) = 87
"001010111",  -- sqrt(7621) = 87
"001010111",  -- sqrt(7622) = 87
"001010111",  -- sqrt(7623) = 87
"001010111",  -- sqrt(7624) = 87
"001010111",  -- sqrt(7625) = 87
"001010111",  -- sqrt(7626) = 87
"001010111",  -- sqrt(7627) = 87
"001010111",  -- sqrt(7628) = 87
"001010111",  -- sqrt(7629) = 87
"001010111",  -- sqrt(7630) = 87
"001010111",  -- sqrt(7631) = 87
"001010111",  -- sqrt(7632) = 87
"001010111",  -- sqrt(7633) = 87
"001010111",  -- sqrt(7634) = 87
"001010111",  -- sqrt(7635) = 87
"001010111",  -- sqrt(7636) = 87
"001010111",  -- sqrt(7637) = 87
"001010111",  -- sqrt(7638) = 87
"001010111",  -- sqrt(7639) = 87
"001010111",  -- sqrt(7640) = 87
"001010111",  -- sqrt(7641) = 87
"001010111",  -- sqrt(7642) = 87
"001010111",  -- sqrt(7643) = 87
"001010111",  -- sqrt(7644) = 87
"001010111",  -- sqrt(7645) = 87
"001010111",  -- sqrt(7646) = 87
"001010111",  -- sqrt(7647) = 87
"001010111",  -- sqrt(7648) = 87
"001010111",  -- sqrt(7649) = 87
"001010111",  -- sqrt(7650) = 87
"001010111",  -- sqrt(7651) = 87
"001010111",  -- sqrt(7652) = 87
"001010111",  -- sqrt(7653) = 87
"001010111",  -- sqrt(7654) = 87
"001010111",  -- sqrt(7655) = 87
"001010111",  -- sqrt(7656) = 87
"001011000",  -- sqrt(7657) = 88
"001011000",  -- sqrt(7658) = 88
"001011000",  -- sqrt(7659) = 88
"001011000",  -- sqrt(7660) = 88
"001011000",  -- sqrt(7661) = 88
"001011000",  -- sqrt(7662) = 88
"001011000",  -- sqrt(7663) = 88
"001011000",  -- sqrt(7664) = 88
"001011000",  -- sqrt(7665) = 88
"001011000",  -- sqrt(7666) = 88
"001011000",  -- sqrt(7667) = 88
"001011000",  -- sqrt(7668) = 88
"001011000",  -- sqrt(7669) = 88
"001011000",  -- sqrt(7670) = 88
"001011000",  -- sqrt(7671) = 88
"001011000",  -- sqrt(7672) = 88
"001011000",  -- sqrt(7673) = 88
"001011000",  -- sqrt(7674) = 88
"001011000",  -- sqrt(7675) = 88
"001011000",  -- sqrt(7676) = 88
"001011000",  -- sqrt(7677) = 88
"001011000",  -- sqrt(7678) = 88
"001011000",  -- sqrt(7679) = 88
"001011000",  -- sqrt(7680) = 88
"001011000",  -- sqrt(7681) = 88
"001011000",  -- sqrt(7682) = 88
"001011000",  -- sqrt(7683) = 88
"001011000",  -- sqrt(7684) = 88
"001011000",  -- sqrt(7685) = 88
"001011000",  -- sqrt(7686) = 88
"001011000",  -- sqrt(7687) = 88
"001011000",  -- sqrt(7688) = 88
"001011000",  -- sqrt(7689) = 88
"001011000",  -- sqrt(7690) = 88
"001011000",  -- sqrt(7691) = 88
"001011000",  -- sqrt(7692) = 88
"001011000",  -- sqrt(7693) = 88
"001011000",  -- sqrt(7694) = 88
"001011000",  -- sqrt(7695) = 88
"001011000",  -- sqrt(7696) = 88
"001011000",  -- sqrt(7697) = 88
"001011000",  -- sqrt(7698) = 88
"001011000",  -- sqrt(7699) = 88
"001011000",  -- sqrt(7700) = 88
"001011000",  -- sqrt(7701) = 88
"001011000",  -- sqrt(7702) = 88
"001011000",  -- sqrt(7703) = 88
"001011000",  -- sqrt(7704) = 88
"001011000",  -- sqrt(7705) = 88
"001011000",  -- sqrt(7706) = 88
"001011000",  -- sqrt(7707) = 88
"001011000",  -- sqrt(7708) = 88
"001011000",  -- sqrt(7709) = 88
"001011000",  -- sqrt(7710) = 88
"001011000",  -- sqrt(7711) = 88
"001011000",  -- sqrt(7712) = 88
"001011000",  -- sqrt(7713) = 88
"001011000",  -- sqrt(7714) = 88
"001011000",  -- sqrt(7715) = 88
"001011000",  -- sqrt(7716) = 88
"001011000",  -- sqrt(7717) = 88
"001011000",  -- sqrt(7718) = 88
"001011000",  -- sqrt(7719) = 88
"001011000",  -- sqrt(7720) = 88
"001011000",  -- sqrt(7721) = 88
"001011000",  -- sqrt(7722) = 88
"001011000",  -- sqrt(7723) = 88
"001011000",  -- sqrt(7724) = 88
"001011000",  -- sqrt(7725) = 88
"001011000",  -- sqrt(7726) = 88
"001011000",  -- sqrt(7727) = 88
"001011000",  -- sqrt(7728) = 88
"001011000",  -- sqrt(7729) = 88
"001011000",  -- sqrt(7730) = 88
"001011000",  -- sqrt(7731) = 88
"001011000",  -- sqrt(7732) = 88
"001011000",  -- sqrt(7733) = 88
"001011000",  -- sqrt(7734) = 88
"001011000",  -- sqrt(7735) = 88
"001011000",  -- sqrt(7736) = 88
"001011000",  -- sqrt(7737) = 88
"001011000",  -- sqrt(7738) = 88
"001011000",  -- sqrt(7739) = 88
"001011000",  -- sqrt(7740) = 88
"001011000",  -- sqrt(7741) = 88
"001011000",  -- sqrt(7742) = 88
"001011000",  -- sqrt(7743) = 88
"001011000",  -- sqrt(7744) = 88
"001011000",  -- sqrt(7745) = 88
"001011000",  -- sqrt(7746) = 88
"001011000",  -- sqrt(7747) = 88
"001011000",  -- sqrt(7748) = 88
"001011000",  -- sqrt(7749) = 88
"001011000",  -- sqrt(7750) = 88
"001011000",  -- sqrt(7751) = 88
"001011000",  -- sqrt(7752) = 88
"001011000",  -- sqrt(7753) = 88
"001011000",  -- sqrt(7754) = 88
"001011000",  -- sqrt(7755) = 88
"001011000",  -- sqrt(7756) = 88
"001011000",  -- sqrt(7757) = 88
"001011000",  -- sqrt(7758) = 88
"001011000",  -- sqrt(7759) = 88
"001011000",  -- sqrt(7760) = 88
"001011000",  -- sqrt(7761) = 88
"001011000",  -- sqrt(7762) = 88
"001011000",  -- sqrt(7763) = 88
"001011000",  -- sqrt(7764) = 88
"001011000",  -- sqrt(7765) = 88
"001011000",  -- sqrt(7766) = 88
"001011000",  -- sqrt(7767) = 88
"001011000",  -- sqrt(7768) = 88
"001011000",  -- sqrt(7769) = 88
"001011000",  -- sqrt(7770) = 88
"001011000",  -- sqrt(7771) = 88
"001011000",  -- sqrt(7772) = 88
"001011000",  -- sqrt(7773) = 88
"001011000",  -- sqrt(7774) = 88
"001011000",  -- sqrt(7775) = 88
"001011000",  -- sqrt(7776) = 88
"001011000",  -- sqrt(7777) = 88
"001011000",  -- sqrt(7778) = 88
"001011000",  -- sqrt(7779) = 88
"001011000",  -- sqrt(7780) = 88
"001011000",  -- sqrt(7781) = 88
"001011000",  -- sqrt(7782) = 88
"001011000",  -- sqrt(7783) = 88
"001011000",  -- sqrt(7784) = 88
"001011000",  -- sqrt(7785) = 88
"001011000",  -- sqrt(7786) = 88
"001011000",  -- sqrt(7787) = 88
"001011000",  -- sqrt(7788) = 88
"001011000",  -- sqrt(7789) = 88
"001011000",  -- sqrt(7790) = 88
"001011000",  -- sqrt(7791) = 88
"001011000",  -- sqrt(7792) = 88
"001011000",  -- sqrt(7793) = 88
"001011000",  -- sqrt(7794) = 88
"001011000",  -- sqrt(7795) = 88
"001011000",  -- sqrt(7796) = 88
"001011000",  -- sqrt(7797) = 88
"001011000",  -- sqrt(7798) = 88
"001011000",  -- sqrt(7799) = 88
"001011000",  -- sqrt(7800) = 88
"001011000",  -- sqrt(7801) = 88
"001011000",  -- sqrt(7802) = 88
"001011000",  -- sqrt(7803) = 88
"001011000",  -- sqrt(7804) = 88
"001011000",  -- sqrt(7805) = 88
"001011000",  -- sqrt(7806) = 88
"001011000",  -- sqrt(7807) = 88
"001011000",  -- sqrt(7808) = 88
"001011000",  -- sqrt(7809) = 88
"001011000",  -- sqrt(7810) = 88
"001011000",  -- sqrt(7811) = 88
"001011000",  -- sqrt(7812) = 88
"001011000",  -- sqrt(7813) = 88
"001011000",  -- sqrt(7814) = 88
"001011000",  -- sqrt(7815) = 88
"001011000",  -- sqrt(7816) = 88
"001011000",  -- sqrt(7817) = 88
"001011000",  -- sqrt(7818) = 88
"001011000",  -- sqrt(7819) = 88
"001011000",  -- sqrt(7820) = 88
"001011000",  -- sqrt(7821) = 88
"001011000",  -- sqrt(7822) = 88
"001011000",  -- sqrt(7823) = 88
"001011000",  -- sqrt(7824) = 88
"001011000",  -- sqrt(7825) = 88
"001011000",  -- sqrt(7826) = 88
"001011000",  -- sqrt(7827) = 88
"001011000",  -- sqrt(7828) = 88
"001011000",  -- sqrt(7829) = 88
"001011000",  -- sqrt(7830) = 88
"001011000",  -- sqrt(7831) = 88
"001011000",  -- sqrt(7832) = 88
"001011001",  -- sqrt(7833) = 89
"001011001",  -- sqrt(7834) = 89
"001011001",  -- sqrt(7835) = 89
"001011001",  -- sqrt(7836) = 89
"001011001",  -- sqrt(7837) = 89
"001011001",  -- sqrt(7838) = 89
"001011001",  -- sqrt(7839) = 89
"001011001",  -- sqrt(7840) = 89
"001011001",  -- sqrt(7841) = 89
"001011001",  -- sqrt(7842) = 89
"001011001",  -- sqrt(7843) = 89
"001011001",  -- sqrt(7844) = 89
"001011001",  -- sqrt(7845) = 89
"001011001",  -- sqrt(7846) = 89
"001011001",  -- sqrt(7847) = 89
"001011001",  -- sqrt(7848) = 89
"001011001",  -- sqrt(7849) = 89
"001011001",  -- sqrt(7850) = 89
"001011001",  -- sqrt(7851) = 89
"001011001",  -- sqrt(7852) = 89
"001011001",  -- sqrt(7853) = 89
"001011001",  -- sqrt(7854) = 89
"001011001",  -- sqrt(7855) = 89
"001011001",  -- sqrt(7856) = 89
"001011001",  -- sqrt(7857) = 89
"001011001",  -- sqrt(7858) = 89
"001011001",  -- sqrt(7859) = 89
"001011001",  -- sqrt(7860) = 89
"001011001",  -- sqrt(7861) = 89
"001011001",  -- sqrt(7862) = 89
"001011001",  -- sqrt(7863) = 89
"001011001",  -- sqrt(7864) = 89
"001011001",  -- sqrt(7865) = 89
"001011001",  -- sqrt(7866) = 89
"001011001",  -- sqrt(7867) = 89
"001011001",  -- sqrt(7868) = 89
"001011001",  -- sqrt(7869) = 89
"001011001",  -- sqrt(7870) = 89
"001011001",  -- sqrt(7871) = 89
"001011001",  -- sqrt(7872) = 89
"001011001",  -- sqrt(7873) = 89
"001011001",  -- sqrt(7874) = 89
"001011001",  -- sqrt(7875) = 89
"001011001",  -- sqrt(7876) = 89
"001011001",  -- sqrt(7877) = 89
"001011001",  -- sqrt(7878) = 89
"001011001",  -- sqrt(7879) = 89
"001011001",  -- sqrt(7880) = 89
"001011001",  -- sqrt(7881) = 89
"001011001",  -- sqrt(7882) = 89
"001011001",  -- sqrt(7883) = 89
"001011001",  -- sqrt(7884) = 89
"001011001",  -- sqrt(7885) = 89
"001011001",  -- sqrt(7886) = 89
"001011001",  -- sqrt(7887) = 89
"001011001",  -- sqrt(7888) = 89
"001011001",  -- sqrt(7889) = 89
"001011001",  -- sqrt(7890) = 89
"001011001",  -- sqrt(7891) = 89
"001011001",  -- sqrt(7892) = 89
"001011001",  -- sqrt(7893) = 89
"001011001",  -- sqrt(7894) = 89
"001011001",  -- sqrt(7895) = 89
"001011001",  -- sqrt(7896) = 89
"001011001",  -- sqrt(7897) = 89
"001011001",  -- sqrt(7898) = 89
"001011001",  -- sqrt(7899) = 89
"001011001",  -- sqrt(7900) = 89
"001011001",  -- sqrt(7901) = 89
"001011001",  -- sqrt(7902) = 89
"001011001",  -- sqrt(7903) = 89
"001011001",  -- sqrt(7904) = 89
"001011001",  -- sqrt(7905) = 89
"001011001",  -- sqrt(7906) = 89
"001011001",  -- sqrt(7907) = 89
"001011001",  -- sqrt(7908) = 89
"001011001",  -- sqrt(7909) = 89
"001011001",  -- sqrt(7910) = 89
"001011001",  -- sqrt(7911) = 89
"001011001",  -- sqrt(7912) = 89
"001011001",  -- sqrt(7913) = 89
"001011001",  -- sqrt(7914) = 89
"001011001",  -- sqrt(7915) = 89
"001011001",  -- sqrt(7916) = 89
"001011001",  -- sqrt(7917) = 89
"001011001",  -- sqrt(7918) = 89
"001011001",  -- sqrt(7919) = 89
"001011001",  -- sqrt(7920) = 89
"001011001",  -- sqrt(7921) = 89
"001011001",  -- sqrt(7922) = 89
"001011001",  -- sqrt(7923) = 89
"001011001",  -- sqrt(7924) = 89
"001011001",  -- sqrt(7925) = 89
"001011001",  -- sqrt(7926) = 89
"001011001",  -- sqrt(7927) = 89
"001011001",  -- sqrt(7928) = 89
"001011001",  -- sqrt(7929) = 89
"001011001",  -- sqrt(7930) = 89
"001011001",  -- sqrt(7931) = 89
"001011001",  -- sqrt(7932) = 89
"001011001",  -- sqrt(7933) = 89
"001011001",  -- sqrt(7934) = 89
"001011001",  -- sqrt(7935) = 89
"001011001",  -- sqrt(7936) = 89
"001011001",  -- sqrt(7937) = 89
"001011001",  -- sqrt(7938) = 89
"001011001",  -- sqrt(7939) = 89
"001011001",  -- sqrt(7940) = 89
"001011001",  -- sqrt(7941) = 89
"001011001",  -- sqrt(7942) = 89
"001011001",  -- sqrt(7943) = 89
"001011001",  -- sqrt(7944) = 89
"001011001",  -- sqrt(7945) = 89
"001011001",  -- sqrt(7946) = 89
"001011001",  -- sqrt(7947) = 89
"001011001",  -- sqrt(7948) = 89
"001011001",  -- sqrt(7949) = 89
"001011001",  -- sqrt(7950) = 89
"001011001",  -- sqrt(7951) = 89
"001011001",  -- sqrt(7952) = 89
"001011001",  -- sqrt(7953) = 89
"001011001",  -- sqrt(7954) = 89
"001011001",  -- sqrt(7955) = 89
"001011001",  -- sqrt(7956) = 89
"001011001",  -- sqrt(7957) = 89
"001011001",  -- sqrt(7958) = 89
"001011001",  -- sqrt(7959) = 89
"001011001",  -- sqrt(7960) = 89
"001011001",  -- sqrt(7961) = 89
"001011001",  -- sqrt(7962) = 89
"001011001",  -- sqrt(7963) = 89
"001011001",  -- sqrt(7964) = 89
"001011001",  -- sqrt(7965) = 89
"001011001",  -- sqrt(7966) = 89
"001011001",  -- sqrt(7967) = 89
"001011001",  -- sqrt(7968) = 89
"001011001",  -- sqrt(7969) = 89
"001011001",  -- sqrt(7970) = 89
"001011001",  -- sqrt(7971) = 89
"001011001",  -- sqrt(7972) = 89
"001011001",  -- sqrt(7973) = 89
"001011001",  -- sqrt(7974) = 89
"001011001",  -- sqrt(7975) = 89
"001011001",  -- sqrt(7976) = 89
"001011001",  -- sqrt(7977) = 89
"001011001",  -- sqrt(7978) = 89
"001011001",  -- sqrt(7979) = 89
"001011001",  -- sqrt(7980) = 89
"001011001",  -- sqrt(7981) = 89
"001011001",  -- sqrt(7982) = 89
"001011001",  -- sqrt(7983) = 89
"001011001",  -- sqrt(7984) = 89
"001011001",  -- sqrt(7985) = 89
"001011001",  -- sqrt(7986) = 89
"001011001",  -- sqrt(7987) = 89
"001011001",  -- sqrt(7988) = 89
"001011001",  -- sqrt(7989) = 89
"001011001",  -- sqrt(7990) = 89
"001011001",  -- sqrt(7991) = 89
"001011001",  -- sqrt(7992) = 89
"001011001",  -- sqrt(7993) = 89
"001011001",  -- sqrt(7994) = 89
"001011001",  -- sqrt(7995) = 89
"001011001",  -- sqrt(7996) = 89
"001011001",  -- sqrt(7997) = 89
"001011001",  -- sqrt(7998) = 89
"001011001",  -- sqrt(7999) = 89
"001011001",  -- sqrt(8000) = 89
"001011001",  -- sqrt(8001) = 89
"001011001",  -- sqrt(8002) = 89
"001011001",  -- sqrt(8003) = 89
"001011001",  -- sqrt(8004) = 89
"001011001",  -- sqrt(8005) = 89
"001011001",  -- sqrt(8006) = 89
"001011001",  -- sqrt(8007) = 89
"001011001",  -- sqrt(8008) = 89
"001011001",  -- sqrt(8009) = 89
"001011001",  -- sqrt(8010) = 89
"001011010",  -- sqrt(8011) = 90
"001011010",  -- sqrt(8012) = 90
"001011010",  -- sqrt(8013) = 90
"001011010",  -- sqrt(8014) = 90
"001011010",  -- sqrt(8015) = 90
"001011010",  -- sqrt(8016) = 90
"001011010",  -- sqrt(8017) = 90
"001011010",  -- sqrt(8018) = 90
"001011010",  -- sqrt(8019) = 90
"001011010",  -- sqrt(8020) = 90
"001011010",  -- sqrt(8021) = 90
"001011010",  -- sqrt(8022) = 90
"001011010",  -- sqrt(8023) = 90
"001011010",  -- sqrt(8024) = 90
"001011010",  -- sqrt(8025) = 90
"001011010",  -- sqrt(8026) = 90
"001011010",  -- sqrt(8027) = 90
"001011010",  -- sqrt(8028) = 90
"001011010",  -- sqrt(8029) = 90
"001011010",  -- sqrt(8030) = 90
"001011010",  -- sqrt(8031) = 90
"001011010",  -- sqrt(8032) = 90
"001011010",  -- sqrt(8033) = 90
"001011010",  -- sqrt(8034) = 90
"001011010",  -- sqrt(8035) = 90
"001011010",  -- sqrt(8036) = 90
"001011010",  -- sqrt(8037) = 90
"001011010",  -- sqrt(8038) = 90
"001011010",  -- sqrt(8039) = 90
"001011010",  -- sqrt(8040) = 90
"001011010",  -- sqrt(8041) = 90
"001011010",  -- sqrt(8042) = 90
"001011010",  -- sqrt(8043) = 90
"001011010",  -- sqrt(8044) = 90
"001011010",  -- sqrt(8045) = 90
"001011010",  -- sqrt(8046) = 90
"001011010",  -- sqrt(8047) = 90
"001011010",  -- sqrt(8048) = 90
"001011010",  -- sqrt(8049) = 90
"001011010",  -- sqrt(8050) = 90
"001011010",  -- sqrt(8051) = 90
"001011010",  -- sqrt(8052) = 90
"001011010",  -- sqrt(8053) = 90
"001011010",  -- sqrt(8054) = 90
"001011010",  -- sqrt(8055) = 90
"001011010",  -- sqrt(8056) = 90
"001011010",  -- sqrt(8057) = 90
"001011010",  -- sqrt(8058) = 90
"001011010",  -- sqrt(8059) = 90
"001011010",  -- sqrt(8060) = 90
"001011010",  -- sqrt(8061) = 90
"001011010",  -- sqrt(8062) = 90
"001011010",  -- sqrt(8063) = 90
"001011010",  -- sqrt(8064) = 90
"001011010",  -- sqrt(8065) = 90
"001011010",  -- sqrt(8066) = 90
"001011010",  -- sqrt(8067) = 90
"001011010",  -- sqrt(8068) = 90
"001011010",  -- sqrt(8069) = 90
"001011010",  -- sqrt(8070) = 90
"001011010",  -- sqrt(8071) = 90
"001011010",  -- sqrt(8072) = 90
"001011010",  -- sqrt(8073) = 90
"001011010",  -- sqrt(8074) = 90
"001011010",  -- sqrt(8075) = 90
"001011010",  -- sqrt(8076) = 90
"001011010",  -- sqrt(8077) = 90
"001011010",  -- sqrt(8078) = 90
"001011010",  -- sqrt(8079) = 90
"001011010",  -- sqrt(8080) = 90
"001011010",  -- sqrt(8081) = 90
"001011010",  -- sqrt(8082) = 90
"001011010",  -- sqrt(8083) = 90
"001011010",  -- sqrt(8084) = 90
"001011010",  -- sqrt(8085) = 90
"001011010",  -- sqrt(8086) = 90
"001011010",  -- sqrt(8087) = 90
"001011010",  -- sqrt(8088) = 90
"001011010",  -- sqrt(8089) = 90
"001011010",  -- sqrt(8090) = 90
"001011010",  -- sqrt(8091) = 90
"001011010",  -- sqrt(8092) = 90
"001011010",  -- sqrt(8093) = 90
"001011010",  -- sqrt(8094) = 90
"001011010",  -- sqrt(8095) = 90
"001011010",  -- sqrt(8096) = 90
"001011010",  -- sqrt(8097) = 90
"001011010",  -- sqrt(8098) = 90
"001011010",  -- sqrt(8099) = 90
"001011010",  -- sqrt(8100) = 90
"001011010",  -- sqrt(8101) = 90
"001011010",  -- sqrt(8102) = 90
"001011010",  -- sqrt(8103) = 90
"001011010",  -- sqrt(8104) = 90
"001011010",  -- sqrt(8105) = 90
"001011010",  -- sqrt(8106) = 90
"001011010",  -- sqrt(8107) = 90
"001011010",  -- sqrt(8108) = 90
"001011010",  -- sqrt(8109) = 90
"001011010",  -- sqrt(8110) = 90
"001011010",  -- sqrt(8111) = 90
"001011010",  -- sqrt(8112) = 90
"001011010",  -- sqrt(8113) = 90
"001011010",  -- sqrt(8114) = 90
"001011010",  -- sqrt(8115) = 90
"001011010",  -- sqrt(8116) = 90
"001011010",  -- sqrt(8117) = 90
"001011010",  -- sqrt(8118) = 90
"001011010",  -- sqrt(8119) = 90
"001011010",  -- sqrt(8120) = 90
"001011010",  -- sqrt(8121) = 90
"001011010",  -- sqrt(8122) = 90
"001011010",  -- sqrt(8123) = 90
"001011010",  -- sqrt(8124) = 90
"001011010",  -- sqrt(8125) = 90
"001011010",  -- sqrt(8126) = 90
"001011010",  -- sqrt(8127) = 90
"001011010",  -- sqrt(8128) = 90
"001011010",  -- sqrt(8129) = 90
"001011010",  -- sqrt(8130) = 90
"001011010",  -- sqrt(8131) = 90
"001011010",  -- sqrt(8132) = 90
"001011010",  -- sqrt(8133) = 90
"001011010",  -- sqrt(8134) = 90
"001011010",  -- sqrt(8135) = 90
"001011010",  -- sqrt(8136) = 90
"001011010",  -- sqrt(8137) = 90
"001011010",  -- sqrt(8138) = 90
"001011010",  -- sqrt(8139) = 90
"001011010",  -- sqrt(8140) = 90
"001011010",  -- sqrt(8141) = 90
"001011010",  -- sqrt(8142) = 90
"001011010",  -- sqrt(8143) = 90
"001011010",  -- sqrt(8144) = 90
"001011010",  -- sqrt(8145) = 90
"001011010",  -- sqrt(8146) = 90
"001011010",  -- sqrt(8147) = 90
"001011010",  -- sqrt(8148) = 90
"001011010",  -- sqrt(8149) = 90
"001011010",  -- sqrt(8150) = 90
"001011010",  -- sqrt(8151) = 90
"001011010",  -- sqrt(8152) = 90
"001011010",  -- sqrt(8153) = 90
"001011010",  -- sqrt(8154) = 90
"001011010",  -- sqrt(8155) = 90
"001011010",  -- sqrt(8156) = 90
"001011010",  -- sqrt(8157) = 90
"001011010",  -- sqrt(8158) = 90
"001011010",  -- sqrt(8159) = 90
"001011010",  -- sqrt(8160) = 90
"001011010",  -- sqrt(8161) = 90
"001011010",  -- sqrt(8162) = 90
"001011010",  -- sqrt(8163) = 90
"001011010",  -- sqrt(8164) = 90
"001011010",  -- sqrt(8165) = 90
"001011010",  -- sqrt(8166) = 90
"001011010",  -- sqrt(8167) = 90
"001011010",  -- sqrt(8168) = 90
"001011010",  -- sqrt(8169) = 90
"001011010",  -- sqrt(8170) = 90
"001011010",  -- sqrt(8171) = 90
"001011010",  -- sqrt(8172) = 90
"001011010",  -- sqrt(8173) = 90
"001011010",  -- sqrt(8174) = 90
"001011010",  -- sqrt(8175) = 90
"001011010",  -- sqrt(8176) = 90
"001011010",  -- sqrt(8177) = 90
"001011010",  -- sqrt(8178) = 90
"001011010",  -- sqrt(8179) = 90
"001011010",  -- sqrt(8180) = 90
"001011010",  -- sqrt(8181) = 90
"001011010",  -- sqrt(8182) = 90
"001011010",  -- sqrt(8183) = 90
"001011010",  -- sqrt(8184) = 90
"001011010",  -- sqrt(8185) = 90
"001011010",  -- sqrt(8186) = 90
"001011010",  -- sqrt(8187) = 90
"001011010",  -- sqrt(8188) = 90
"001011010",  -- sqrt(8189) = 90
"001011010",  -- sqrt(8190) = 90
"001011011"  -- sqrt(8191) = 91
    );

begin
    process(Clk)
    begin
        if rising_edge(Clk) then
            if en = '1' then
                --take the last 13 bits because it seems like VHD files have a 10000 line limit
                SqRoot <= ROM(to_integer(unsigned(Addr(12 downto 0))));
                data_valid <= '1';
            else
                data_valid <= '0';
            end if;
        end if;
    end process;
end architecture;
